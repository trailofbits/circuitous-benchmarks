module circuit(
input [1854:0] current,
input [1854:0] next,

output [0:0] result,
output [0:0] dummy
);
wire [31:0] Advice_1 = current[31: 0];
wire [2:0] Advice_10 = current[34: 32];
wire [2:0] Advice_11 = current[37: 35];
wire [2:0] Advice_12 = current[40: 38];
wire [2:0] Advice_13 = current[43: 41];
wire [1:0] Advice_14 = current[45: 44];
wire [1:0] Advice_15 = current[47: 46];
wire [2:0] Advice_16 = current[50: 48];
wire Advice_17 = current[51: 51];
wire [2:0] Advice_18 = current[54: 52];
wire Advice_19 = current[55: 55];
wire [63:0] Advice_2 = current[119: 56];
wire Advice_20 = current[120: 120];
wire Advice_21 = current[121: 121];
wire [1:0] Advice_22 = current[123: 122];
wire [1:0] Advice_23 = current[125: 124];
wire [2:0] Advice_24 = current[128: 126];
wire [1:0] Advice_25 = current[130: 129];
wire Advice_26 = current[131: 131];
wire [2:0] Advice_27 = current[134: 132];
wire [2:0] Advice_28 = current[137: 135];
wire [2:0] Advice_29 = current[140: 138];
wire [63:0] Advice_3 = current[204: 141];
wire [2:0] Advice_30 = current[207: 205];
wire [2:0] Advice_31 = current[210: 208];
wire Advice_32 = current[211: 211];
wire [1:0] Advice_33 = current[213: 212];
wire Advice_34 = current[214: 214];
wire [2:0] Advice_4 = current[217: 215];
wire [2:0] Advice_5 = current[220: 218];
wire [31:0] Advice_6 = current[252: 221];
wire [2:0] Advice_7 = current[255: 253];
wire [2:0] Advice_8 = current[258: 256];
wire [31:0] Advice_9 = current[290: 259];
wire In_error_flag = current[291: 291];
wire In_register_AF = current[620: 620];
wire [31:0] In_register_CSBASE = current[653: 622];
wire [7:0] In_register_DF = current[661: 654];
wire [31:0] In_register_DSBASE = current[693: 662];
wire [31:0] In_register_EAX = current[725: 694];
wire [31:0] In_register_EBP = current[757: 726];
wire [31:0] In_register_EBX = current[789: 758];
wire [31:0] In_register_ECX = current[821: 790];
wire [31:0] In_register_EDI = current[853: 822];
wire [31:0] In_register_EDX = current[885: 854];
wire [31:0] In_register_EIP = current[917: 886];
wire [31:0] In_register_ESBASE = current[949: 918];
wire [31:0] In_register_ESI = current[981: 950];
wire [31:0] In_register_ESP = current[1013: 982];
wire [31:0] In_register_FSBASE = current[1045: 1014];
wire [31:0] In_register_GSBASE = current[1077: 1046];
wire In_register_PF = current[1079: 1079];
wire In_register_SF = current[1080: 1080];
wire [31:0] In_register_SSBASE = current[1112: 1081];
wire In_register_ZF = current[1113: 1113];
wire [63:0] In_timestamp = current[1177: 1114];
wire Out_error_flag = next[291: 291];
wire Out_register_AF = next[620: 620];
wire Out_register_CF = next[621: 621];
wire [31:0] Out_register_CSBASE = next[653: 622];
wire [7:0] Out_register_DF = next[661: 654];
wire [31:0] Out_register_DSBASE = next[693: 662];
wire [31:0] Out_register_EAX = next[725: 694];
wire [31:0] Out_register_EBP = next[757: 726];
wire [31:0] Out_register_EBX = next[789: 758];
wire [31:0] Out_register_ECX = next[821: 790];
wire [31:0] Out_register_EDI = next[853: 822];
wire [31:0] Out_register_EDX = next[885: 854];
wire [31:0] Out_register_EIP = next[917: 886];
wire [31:0] Out_register_ESBASE = next[949: 918];
wire [31:0] Out_register_ESI = next[981: 950];
wire [31:0] Out_register_ESP = next[1013: 982];
wire [31:0] Out_register_FSBASE = next[1045: 1014];
wire [31:0] Out_register_GSBASE = next[1077: 1046];
wire Out_register_OF = next[1078: 1078];
wire Out_register_PF = next[1079: 1079];
wire Out_register_SF = next[1080: 1080];
wire [31:0] Out_register_SSBASE = next[1112: 1081];
wire Out_register_ZF = next[1113: 1113];
wire [63:0] Out_timestamp = next[1177: 1114];
wire [119:0] instruction_bits = current[411: 292];
wire [207:0] memory_0 = current[619: 412];
wire [31:0] v4 = 32'b00000000000000000000000000000000;
wire [31:0] v6 = In_register_DSBASE + v4;
wire [31:0] v7 = v4 << v4;
wire [31:0] v8 = v6 + v7;
wire [31:0] va = instruction_bits[63: 32];
wire [31:0] vc = v8 + va;
wire ve = vc == Advice_1;
wire vf = 1'b0;
wire v11 = vf == Out_error_flag;
wire v13 = In_error_flag == vf;
wire [31:0] v15 = 32'b00000000000000001111111111111111;
wire [31:0] v16 = In_register_EAX & v15;
wire [63:0] v19 = Advice_2 * Advice_3;
wire [31:0] v1a = v19[31:0];
wire [15:0] v1b = v1a[15:0];
wire [31:0] v1c = { 16'b0000000000000000, v1b };
wire [31:0] v1d = v16 | v1c;
wire v1f = v1d == Out_register_EAX;
wire v22 = In_register_EBX == Out_register_EBX;
wire v25 = In_register_ECX == Out_register_ECX;
wire [31:0] v27 = In_register_EDX & v15;
wire [31:0] v28 = 32'b00001000000000000000000000000000;
wire [31:0] v29 = v1a >> v28;
wire [15:0] v2a = v29[15:0];
wire [31:0] v2b = { 16'b0000000000000000, v2a };
wire [31:0] v2c = v27 | v2b;
wire v2e = v2c == Out_register_EDX;
wire v31 = In_register_ESI == Out_register_ESI;
wire v34 = In_register_EDI == Out_register_EDI;
wire v37 = In_register_ESP == Out_register_ESP;
wire v3a = In_register_EBP == Out_register_EBP;
wire [31:0] v3c = 32'b00010000000000000000000000000000;
wire [31:0] v3d = In_register_EIP + v3c;
wire v3f = v3d == Out_register_EIP;
wire v42 = In_register_CSBASE == Out_register_CSBASE;
wire v45 = In_register_SSBASE == Out_register_SSBASE;
wire v48 = In_register_ESBASE == Out_register_ESBASE;
wire v4a = In_register_DSBASE == Out_register_DSBASE;
wire v4d = In_register_GSBASE == Out_register_GSBASE;
wire v50 = In_register_FSBASE == Out_register_FSBASE;
wire v53 = In_register_AF == Out_register_AF;
wire [31:0] v54 = 32'b00000000000000011111111111111111;
wire [31:0] v55 = v1a + v54;
wire v56 = v55 < v15;
wire v58 = v56 == Out_register_CF;
wire v5b = In_register_DF == Out_register_DF;
wire v5d = v56 == Out_register_OF;
wire v60 = In_register_PF == Out_register_PF;
wire v63 = In_register_SF == Out_register_SF;
wire v66 = In_register_ZF == Out_register_ZF;
wire v67 = v1f & v22 & v25 & v2e & v31 & v34 & v37 & v3a & v3f & v42 & v45 & v48 & v4a & v4d & v50 & v53 & v58 & v5b & v5d & v60 & v63 & v66;
wire [3:0] v69 = 4'b0100;
wire v6b =  v69 == memory_0[15: 12] && Advice_1 == memory_0[79: 16] && In_timestamp == memory_0[207: 144] && 4'd0 == memory_0[11: 8] && 1'b1 == memory_0[0: 0] && 6'b000000 == memory_0[7: 2] && 1'b0 == memory_0[1: 1];
wire [31:0] v6c = 32'b01100110011001101110111110110100;
wire [31:0] v6d = instruction_bits[31: 0];
wire v6e = v6c == v6d;
wire [55:0] v6f = 56'b00000000000000000000000000000000000000000000000000000000;
wire [55:0] v70 = instruction_bits[119: 64];
wire v71 = v6f == v70;
wire v72 = 1'b1;
wire v73 = v72 & v72 & v72;
wire v74 = v6e & v71 & v73;
wire [63:0] v75 = 64'b1000000000000000000000000000000000000000000000000000000000000000;
wire [63:0] v76 = In_timestamp + v75;
wire v78 = v76 == Out_timestamp;
wire v79 = In_error_flag ^ v72;
wire v7a = v79 | Out_error_flag;
wire [31:0] v7b = memory_0[79: 48];
wire [15:0] v7c = v7b[15:0];
wire [15:0] pad_125 = (v7c[15:15] == 1'b1) ?16'b1111111111111111 : 16'b0000000000000000;
wire [31:0] v7d = { pad_125, v7c };
wire [31:0] pad_126 = (v7d[31:31] == 1'b1) ?32'b11111111111111111111111111111111 : 32'b00000000000000000000000000000000;
wire [63:0] v7e = { pad_126, v7d };
wire v7f = v7e == Advice_2;
wire [15:0] v80 = In_register_EAX[15:0];
wire [15:0] pad_129 = (v80[15:15] == 1'b1) ?16'b1111111111111111 : 16'b0000000000000000;
wire [31:0] v81 = { pad_129, v80 };
wire [31:0] pad_130 = (v81[31:31] == 1'b1) ?32'b11111111111111111111111111111111 : 32'b00000000000000000000000000000000;
wire [63:0] v82 = { pad_130, v81 };
wire v83 = v82 == Advice_3;
wire v84 = ve & v11 & v13 & v67 & v6b & v74 & v78 & v7a & v7f & v83;
wire rnx2x0 = 1'b0 || v84;
wire onx2x0 = 1'b0 || ( 1'b0 && v84);
wire [31:0] v85 = instruction_bits[47: 16];
wire [31:0] v87 = v8 + v85;
wire v88 = v87 == Advice_1;
wire [3:0] v89 = 4'b0010;
wire v8a =  v89 == memory_0[15: 12] && Advice_1 == memory_0[79: 16] && In_timestamp == memory_0[207: 144] && 4'd0 == memory_0[11: 8] && 1'b1 == memory_0[0: 0] && 6'b000000 == memory_0[7: 2] && 1'b0 == memory_0[1: 1];
wire v8b = v1a == Out_register_EAX;
wire [63:0] v8c = 64'b0000010000000000000000000000000000000000000000000000000000000000;
wire [63:0] v8d = v19 >> v8c;
wire [31:0] v8e = v8d[31:0];
wire v8f = v8e == Out_register_EDX;
wire [31:0] v90 = 32'b01100000000000000000000000000000;
wire [31:0] v91 = In_register_EIP + v90;
wire v92 = v91 == Out_register_EIP;
wire [63:0] v93 = 64'b0000000000000000000000000000000111111111111111111111111111111111;
wire [63:0] v94 = v19 + v93;
wire [63:0] v95 = 64'b0000000000000000000000000000000011111111111111111111111111111111;
wire v96 = v94 < v95;
wire v97 = v96 == Out_register_CF;
wire v98 = v96 == Out_register_OF;
wire v99 = v8b & v22 & v25 & v8f & v31 & v34 & v37 & v3a & v92 & v42 & v45 & v48 & v4a & v4d & v50 & v53 & v97 & v5b & v98 & v60 & v63 & v66;
wire [15:0] v9a = 16'b1110111110110100;
wire [15:0] v9b = instruction_bits[15: 0];
wire v9c = v9a == v9b;
wire [71:0] v9d = 72'b000000000000000000000000000000000000000000000000000000000000000000000000;
wire [71:0] v9e = instruction_bits[119: 48];
wire v9f = v9d == v9e;
wire va0 = v9c & v9f & v73;
wire [31:0] pad_161 = (v7b[31:31] == 1'b1) ?32'b11111111111111111111111111111111 : 32'b00000000000000000000000000000000;
wire [63:0] va1 = { pad_161, v7b };
wire va2 = va1 == Advice_2;
wire [31:0] pad_163 = (In_register_EAX[31:31] == 1'b1) ?32'b11111111111111111111111111111111 : 32'b00000000000000000000000000000000;
wire [63:0] va3 = { pad_163, In_register_EAX };
wire va4 = va3 == Advice_3;
wire va5 = v88 & v11 & v8a & v13 & v99 & va0 & v78 & v7a & va2 & va4;
wire rnx2x1 = rnx2x0 || va5;
wire onx2x1 = onx2x0 || ( rnx2x0 && va5);
wire [31:0] va6 = instruction_bits[55: 24];
wire [31:0] va8 = v8 + va6;
wire va9 = va8 == Advice_1;
wire [31:0] vaa = 32'b11100000000000000000000000000000;
wire [31:0] vab = In_register_EIP + vaa;
wire vac = vab == Out_register_EIP;
wire vad = v8b & v22 & v25 & v8f & v31 & v34 & v37 & v3a & vac & v42 & v45 & v48 & v4a & v4d & v50 & v53 & v97 & v5b & v98 & v60 & v63 & v66;
wire [23:0] vae = 24'b111011110011010010100110;
wire [23:0] vaf = instruction_bits[23: 0];
wire vb0 = vae == vaf;
wire [63:0] vb1 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
wire [63:0] vb2 = instruction_bits[119: 56];
wire vb3 = vb1 == vb2;
wire vb4 = vb0 & vb3 & v73;
wire vb5 = va9 & vad & v13 & v8a & v78 & v11 & vb4 & v7a & va2 & va4;
wire rnx2x2 = rnx2x1 || vb5;
wire onx2x2 = onx2x1 || ( rnx2x1 && vb5);
wire [31:0] vb6 = 32'b00000000111111111111111111111111;
wire [31:0] vb7 = In_register_EAX & vb6;
wire [15:0] vb8 = v19[15:0];
wire [7:0] vb9 = vb8[7:0];
wire [31:0] vba = { 24'b000000000000000000000000, vb9 };
wire [31:0] vbb = vb7 | vba;
wire [31:0] vbc = 32'b11111111000000001111111111111111;
wire [31:0] vbd = vbb & vbc;
wire [15:0] vbe = 16'b0001000000000000;
wire [15:0] vbf = vb8 >> vbe;
wire [7:0] vc0 = vbf[7:0];
wire [31:0] vc1 = { 24'b000000000000000000000000, vc0 };
wire [31:0] vc2 = vc1 << v3c;
wire [31:0] vc3 = vbd | vc2;
wire vc4 = vc3 == Out_register_EAX;
wire vc5 = In_register_EDX == Out_register_EDX;
wire [15:0] vc6 = 16'b1111111100000000;
wire vc7 = vb8 > vc6;
wire vc8 = vc7 == Out_register_CF;
wire vc9 = vc7 == Out_register_OF;
wire vca = vc4 & v22 & v25 & vc5 & v31 & v34 & v37 & v3a & v92 & v42 & v45 & v48 & v4a & v4d & v50 & v53 & vc8 & v5b & vc9 & v60 & v63 & v66;
wire [15:0] vcb = 16'b0110111110100100;
wire vcc = vcb == v9b;
wire vcd = vcc & v9f & v73;
wire [3:0] vce = 4'b1000;
wire vcf =  vce == memory_0[15: 12] && Advice_1 == memory_0[79: 16] && In_timestamp == memory_0[207: 144] && 4'd0 == memory_0[11: 8] && 1'b1 == memory_0[0: 0] && 6'b000000 == memory_0[7: 2] && 1'b0 == memory_0[1: 1];
wire [7:0] vd0 = v7b[7:0];
wire [15:0] vd1 = { 8'b00000000, vd0 };
wire [15:0] pad_210 = (vd1[15:15] == 1'b1) ?48'b111111111111111111111111111111111111111111111111 : 48'b000000000000000000000000000000000000000000000000;
wire [63:0] vd2 = { pad_210, vd1 };
wire vd3 = vd2 == Advice_2;
wire [7:0] vd4 = In_register_EAX[7:0];
wire [15:0] vd5 = { 8'b00000000, vd4 };
wire [15:0] pad_214 = (vd5[15:15] == 1'b1) ?48'b111111111111111111111111111111111111111111111111 : 48'b000000000000000000000000000000000000000000000000;
wire [63:0] vd6 = { pad_214, vd5 };
wire vd7 = vd6 == Advice_3;
wire vd8 = v88 & vca & v11 & v13 & vcd & vcf & v78 & v7a & vd3 & vd7;
wire rnx2x3 = rnx2x2 || vd8;
wire onx2x3 = onx2x2 || ( rnx2x2 && vd8);
wire [31:0] vd9 = 32'b00100000000000000000000000000000;
wire [31:0] vda = In_register_EIP + vd9;
wire vdb = vda == Out_register_EIP;
wire vdc = v1f & v22 & v25 & v2e & v31 & v34 & v37 & v3a & vdb & v42 & v45 & v48 & v4a & v4d & v50 & v53 & v58 & v5b & v5d & v60 & v63 & v66;
wire [2:0] vdd = instruction_bits[26: 24];
wire [2:0] vde = { vdd };
wire ve0 = vde == Advice_4;
wire [31:0] ve2 = ( Advice_5 == 3'd0) ? In_register_EAX :
	( Advice_5 == 3'd1) ? In_register_ECX :
	( Advice_5 == 3'd2) ? In_register_EDX :
	( Advice_5 == 3'd3) ? In_register_EBX :
	( Advice_5 == 3'd4) ? In_register_ESP :
	( Advice_5 == 3'd5) ? In_register_EBP :
	( Advice_5 == 3'd6) ? In_register_ESI : In_register_EDI;
wire [31:0] ve3 = 32'b11111111111111110000000000000000;
wire [31:0] ve4 = ve2 & ve3;
wire ve5 = ve4 == Advice_1;
wire [23:0] ve6 = 24'b011001100110011011101111;
wire ve7 = ve6 == vaf;
wire [4:0] ve8 = 5'b10111;
wire [4:0] ve9 = instruction_bits[31: 27];
wire vea = ve8 == ve9;
wire [87:0] veb = 88'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
wire [87:0] vec = instruction_bits[119: 32];
wire ved = veb == vec;
wire vee = v72;
wire vef = ve7 & vea & ved & vee;
wire vf0 = Advice_4 == Advice_5;
wire [31:0] vf1 = Advice_1 << v28;
wire [31:0] vf2 = vf1 >>> v28;
wire [31:0] pad_243 = (vf2[31:31] == 1'b1) ?32'b11111111111111111111111111111111 : 32'b00000000000000000000000000000000;
wire [63:0] vf3 = { pad_243, vf2 };
wire vf4 = vf3 == Advice_2;
wire vf5 = v11 & vdc & v13 & v7a & ve0 & ve5 & vef & v78 & vf0 & vf4 & v83;
wire rnx2x4 = rnx2x3 || vf5;
wire onx2x4 = onx2x3 || ( rnx2x3 && vf5);
wire [31:0] vf6 = 32'b01000000000000000000000000000000;
wire [31:0] vf7 = In_register_EIP + vf6;
wire vf8 = vf7 == Out_register_EIP;
wire vf9 = v8b & v22 & v25 & v8f & v31 & v34 & v37 & v3a & vf8 & v42 & v45 & v48 & v4a & v4d & v50 & v53 & v97 & v5b & v98 & v60 & v63 & v66;
wire vfa = ve2 == Advice_1;
wire [2:0] vfb = instruction_bits[10: 8];
wire [2:0] vfc = { vfb };
wire vfd = vfc == Advice_4;
wire [7:0] vfe = 8'b11101111;
wire [7:0] vff = instruction_bits[7: 0];
wire v100 = vfe == vff;
wire [4:0] v101 = instruction_bits[15: 11];
wire v102 = ve8 == v101;
wire [103:0] v103 = 104'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
wire [103:0] v104 = instruction_bits[119: 16];
wire v105 = v103 == v104;
wire v106 = v100 & v102 & v105 & vee;
wire v107 = va3 == Advice_2;
wire [31:0] pad_264 = (Advice_1[31:31] == 1'b1) ?32'b11111111111111111111111111111111 : 32'b00000000000000000000000000000000;
wire [63:0] v108 = { pad_264, Advice_1 };
wire v109 = v108 == Advice_3;
wire v10a = vf9 & vfa & v11 & v13 & v7a & vfd & v106 & v78 & vf0 & v107 & v109;
wire rnx2x5 = rnx2x4 || v10a;
wire onx2x5 = onx2x4 || ( rnx2x4 && v10a);
wire [31:0] v10b = 32'b11000000000000000000000000000000;
wire [31:0] v10c = In_register_EIP + v10b;
wire v10d = v10c == Out_register_EIP;
wire v10e = v8b & v22 & v25 & v8f & v31 & v34 & v37 & v3a & v10d & v42 & v45 & v48 & v4a & v4d & v50 & v53 & v97 & v5b & v98 & v60 & v63 & v66;
wire [15:0] v10f = 16'b1110011011101111;
wire v110 = v10f == v9b;
wire [4:0] v111 = instruction_bits[23: 19];
wire v112 = ve8 == v111;
wire [95:0] v113 = 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
wire [95:0] v114 = instruction_bits[119: 24];
wire v115 = v113 == v114;
wire v116 = v110 & v112 & v115 & vee;
wire [2:0] v117 = instruction_bits[18: 16];
wire [2:0] v118 = { v117 };
wire v119 = v118 == Advice_4;
wire v11a = v10e & vfa & v13 & v116 & v11 & v119 & v78 & v7a & vf0 & v107 & v109;
wire rnx2x6 = rnx2x5 || v11a;
wire onx2x6 = onx2x5 || ( rnx2x5 && v11a);
wire [7:0] v11b = instruction_bits[23: 16];
wire [7:0] pad_284 = (v11b[7:7] == 1'b1) ?24'b111111111111111111111111 : 24'b000000000000000000000000;
wire [31:0] v11c = { pad_284, v11b };
wire v11f = v11c == Advice_6;
wire [7:0] v120 = 8'b11010110;
wire v121 = v120 == vff;
wire [1:0] v122 = 2'b11;
wire [1:0] v123 = instruction_bits[15: 14];
wire v124 = v122 == v123;
wire v125 = v121 & v124 & v115 & v72;
wire v127 = vfc == Advice_7;
wire [31:0] v128 = { v1a };
wire [31:0] v12a = ( Advice_8 == 3'd0) ? Out_register_EAX :
	( Advice_8 == 3'd1) ? Out_register_ECX :
	( Advice_8 == 3'd2) ? Out_register_EDX :
	( Advice_8 == 3'd3) ? Out_register_EBX :
	( Advice_8 == 3'd4) ? Out_register_ESP :
	( Advice_8 == 3'd5) ? Out_register_EBP :
	( Advice_8 == 3'd6) ? Out_register_ESI : Out_register_EDI;
wire v12b = v128 == v12a;
wire [2:0] v12c = 3'b000;
wire v12d = Advice_4 == v12c;
wire v12e = In_register_EAX == Out_register_EAX;
wire v12f = v12d | v12e;
wire [2:0] v130 = 3'b110;
wire v131 = Advice_4 == v130;
wire v132 = v131 | v22;
wire [2:0] v133 = 3'b100;
wire v134 = Advice_4 == v133;
wire v135 = v134 | v25;
wire [2:0] v136 = 3'b010;
wire v137 = Advice_4 == v136;
wire v138 = v137 | vc5;
wire [2:0] v139 = 3'b011;
wire v13a = Advice_4 == v139;
wire v13b = v13a | v31;
wire [2:0] v13c = 3'b111;
wire v13d = Advice_4 == v13c;
wire v13e = v13d | v34;
wire [2:0] v13f = 3'b001;
wire v140 = Advice_4 == v13f;
wire v141 = v140 | v37;
wire [2:0] v142 = 3'b101;
wire v143 = Advice_4 == v142;
wire v144 = v143 | v3a;
wire v145 = v12f & v132 & v135 & v138 & v13b & v13e & v141 & v144 & v10d & v42 & v45 & v48 & v4a & v4d & v50 & v53 & v97 & v5b & v98 & v60 & v63 & v66;
wire v146 = v12b & v145;
wire v148 = ve2 == Advice_9;
wire [2:0] v149 = instruction_bits[13: 11];
wire [2:0] v14a = { v149 };
wire v14b = v14a == Advice_4;
wire v14c = Advice_7 == Advice_5;
wire v14d = Advice_4 == Advice_8;
wire [31:0] pad_334 = (Advice_6[31:31] == 1'b1) ?32'b11111111111111111111111111111111 : 32'b00000000000000000000000000000000;
wire [63:0] v14e = { pad_334, Advice_6 };
wire v14f = v14e == Advice_2;
wire [31:0] pad_336 = (Advice_9[31:31] == 1'b1) ?32'b11111111111111111111111111111111 : 32'b00000000000000000000000000000000;
wire [63:0] v150 = { pad_336, Advice_9 };
wire v151 = v150 == Advice_3;
wire v152 = v11f & v13 & v125 & v127 & v146 & v78 & v148 & v11 & v14b & v7a & v14c & v14d & v14f & v151;
wire rnx2x7 = rnx2x6 || v152;
wire onx2x7 = onx2x6 || ( rnx2x6 && v152);
wire v153 = v12f & v132 & v135 & v138 & v13b & v13e & v141 & v144 & vdb & v42 & v45 & v48 & v4a & v4d & v50 & v53 & v97 & v5b & v98 & v60 & v63 & v66;
wire v154 = v12b & v153;
wire [7:0] v155 = instruction_bits[31: 24];
wire [7:0] pad_342 = (v155[7:7] == 1'b1) ?24'b111111111111111111111111 : 24'b000000000000000000000000;
wire [31:0] v156 = { pad_342, v155 };
wire v158 = v156 == Advice_6;
wire v159 = v118 == Advice_7;
wire [2:0] v15a = instruction_bits[21: 19];
wire [2:0] v15b = { v15a };
wire v15c = v15b == Advice_4;
wire [15:0] v15d = 16'b0110010011010110;
wire v15e = v15d == v9b;
wire [1:0] v15f = instruction_bits[23: 22];
wire v160 = v122 == v15f;
wire v161 = v15e & v160 & ved & v72;
wire v162 = v154 & v148 & v11 & v158 & v159 & v15c & v161 & v13 & v78 & v7a & v14c & v14d & v14f & v151;
wire rnx2x8 = rnx2x7 || v162;
wire onx2x8 = onx2x7 || ( rnx2x7 && v162);
wire [2:0] v163 = instruction_bits[29: 27];
wire [2:0] v164 = { v163 };
wire v165 = v164 == Advice_4;
wire [23:0] v166 = 24'b101001101110011011010110;
wire v167 = v166 == vaf;
wire [1:0] v168 = instruction_bits[31: 30];
wire v169 = v122 == v168;
wire [79:0] v16a = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
wire [79:0] v16b = instruction_bits[119: 40];
wire v16c = v16a == v16b;
wire v16d = v167 & v169 & v16c & v72;
wire [31:0] v16e = 32'b10100000000000000000000000000000;
wire [31:0] v16f = In_register_EIP + v16e;
wire v170 = v16f == Out_register_EIP;
wire v171 = v12f & v132 & v135 & v138 & v13b & v13e & v141 & v144 & v170 & v42 & v45 & v48 & v4a & v4d & v50 & v53 & v97 & v5b & v98 & v60 & v63 & v66;
wire v172 = v12b & v171;
wire [7:0] v173 = instruction_bits[39: 32];
wire [7:0] pad_372 = (v173[7:7] == 1'b1) ?24'b111111111111111111111111 : 24'b000000000000000000000000;
wire [31:0] v174 = { pad_372, v173 };
wire v176 = v174 == Advice_6;
wire v177 = vde == Advice_7;
wire v178 = v11 & v148 & v13 & v165 & v16d & v172 & v78 & v176 & v177 & v7a & v14c & v14d & v14f & v151;
wire rnx2x9 = rnx2x8 || v178;
wire onx2x9 = onx2x8 || ( rnx2x8 && v178);
wire [15:0] v179 = instruction_bits[39: 24];
wire [15:0] pad_378 = (v179[15:15] == 1'b1) ?16'b1111111111111111 : 16'b0000000000000000;
wire [31:0] v17a = { pad_378, v179 };
wire v17c = v17a == Advice_6;
wire v17d = ve4 == Advice_9;
wire [31:0] v17f = ( Advice_10 == 3'd0) ? In_register_EAX :
	( Advice_10 == 3'd1) ? In_register_ECX :
	( Advice_10 == 3'd2) ? In_register_EDX :
	( Advice_10 == 3'd3) ? In_register_EBX :
	( Advice_10 == 3'd4) ? In_register_ESP :
	( Advice_10 == 3'd5) ? In_register_EBP :
	( Advice_10 == 3'd6) ? In_register_ESI : In_register_EDI;
wire [15:0] v180 = v17f[31: 16];
wire [31:0] v181 = { v180 , v1b };
wire v182 = v181 == v12a;
wire v183 = v12f & v132 & v135 & v138 & v13b & v13e & v141 & v144 & v170 & v42 & v45 & v48 & v4a & v4d & v50 & v53 & v58 & v5b & v5d & v60 & v63 & v66;
wire v184 = v182 & v183;
wire [15:0] v185 = 16'b0110011010010110;
wire v186 = v185 == v9b;
wire v187 = v186 & v160 & v16c & v72;
wire v188 = Advice_4 == Advice_10;
wire [31:0] v189 = Advice_6 << v28;
wire [31:0] v18a = v189 >>> v28;
wire [31:0] pad_395 = (v18a[31:31] == 1'b1) ?32'b11111111111111111111111111111111 : 32'b00000000000000000000000000000000;
wire [63:0] v18b = { pad_395, v18a };
wire v18c = v18b == Advice_2;
wire [31:0] v18d = Advice_9 << v28;
wire [31:0] v18e = v18d >>> v28;
wire [31:0] pad_399 = (v18e[31:31] == 1'b1) ?32'b11111111111111111111111111111111 : 32'b00000000000000000000000000000000;
wire [63:0] v18f = { pad_399, v18e };
wire v190 = v18f == Advice_3;
wire v191 = v17c & v17d & v11 & v184 & v13 & v15c & v78 & v159 & v187 & v7a & v14c & v188 & v14d & v18c & v190;
wire rnx2x10 = rnx2x9 || v191;
wire onx2x10 = onx2x9 || ( rnx2x9 && v191);
wire v192 = v12f & v132 & v135 & v138 & v13b & v13e & v141 & v144 & v92 & v42 & v45 & v48 & v4a & v4d & v50 & v53 & v58 & v5b & v5d & v60 & v63 & v66;
wire v193 = v182 & v192;
wire [23:0] v194 = 24'b011001000110011010010110;
wire v195 = v194 == vaf;
wire v196 = v195 & v169 & v9f & v72;
wire [15:0] v197 = instruction_bits[47: 32];
wire [15:0] pad_408 = (v197[15:15] == 1'b1) ?16'b1111111111111111 : 16'b0000000000000000;
wire [31:0] v198 = { pad_408, v197 };
wire v19a = v198 == Advice_6;
wire v19b = v193 & v196 & v19a & v17d & v78 & v177 & v165 & v11 & v13 & v7a & v14c & v14d & v188 & v18c & v190;
wire rnx2x11 = rnx2x10 || v19b;
wire onx2x11 = onx2x10 || ( rnx2x10 && v19b);
wire v19c = v85 == Advice_6;
wire v19d = v12f & v132 & v135 & v138 & v13b & v13e & v141 & v144 & v92 & v42 & v45 & v48 & v4a & v4d & v50 & v53 & v97 & v5b & v98 & v60 & v63 & v66;
wire v19e = v12b & v19d;
wire [7:0] v19f = 8'b10010110;
wire v1a0 = v19f == vff;
wire v1a1 = v1a0 & v124 & v9f & v72;
wire v1a2 = v19c & v148 & v11 & v13 & v14b & v127 & v19e & v1a1 & v78 & v7a & v14c & v14d & v14f & v151;
wire rnx2x12 = rnx2x11 || v1a2;
wire onx2x12 = onx2x11 || ( rnx2x11 && v1a2);
wire v1a3 = v12f & v132 & v135 & v138 & v13b & v13e & v141 & v144 & vac & v42 & v45 & v48 & v4a & v4d & v50 & v53 & v97 & v5b & v98 & v60 & v63 & v66;
wire v1a4 = v12b & v1a3;
wire v1a5 = va6 == Advice_6;
wire [15:0] v1a6 = 16'b1110011010010110;
wire v1a7 = v1a6 == v9b;
wire v1a8 = v1a7 & v160 & vb3 & v72;
wire v1a9 = v1a4 & v1a5 & v148 & v1a8 & v159 & v78 & v11 & v13 & v15c & v7a & v14c & v14d & v14f & v151;
wire rnx2x13 = rnx2x12 || v1a9;
wire onx2x13 = onx2x12 || ( rnx2x12 && v1a9);
wire v1aa = va == Advice_6;
wire [23:0] v1ab = 24'b101001100010011010010110;
wire v1ac = v1ab == vaf;
wire v1ad = v1ac & v169 & v71 & v72;
wire v1ae = v12f & v132 & v135 & v138 & v13b & v13e & v141 & v144 & v3f & v42 & v45 & v48 & v4a & v4d & v50 & v53 & v97 & v5b & v98 & v60 & v63 & v66;
wire v1af = v12b & v1ae;
wire v1b0 = v148 & v11 & v1aa & v13 & v177 & v165 & v1ad & v78 & v1af & v7a & v14c & v14d & v14f & v151;
wire rnx2x14 = rnx2x13 || v1b0;
wire onx2x14 = onx2x13 || ( rnx2x13 && v1b0);
wire [31:0] v1b2 = ( Advice_11 == 3'd0) ? In_register_DSBASE :
	( Advice_11 == 3'd1) ? In_register_DSBASE :
	( Advice_11 == 3'd2) ? In_register_DSBASE :
	( Advice_11 == 3'd3) ? In_register_DSBASE :
	( Advice_11 == 3'd4) ? In_register_SSBASE :
	( Advice_11 == 3'd5) ? In_register_SSBASE :
	( Advice_11 == 3'd6) ? In_register_DSBASE : In_register_DSBASE;
wire [31:0] v1b3 = v1b2 + ve2;
wire [31:0] v1b4 = v1b3 + v7;
wire [31:0] v1b5 = v1b4 + v4;
wire v1b6 = v1b5 == Advice_9;
wire v1b8 = vfc == Advice_12;
wire v1b9 =  v89 == memory_0[15: 12] && Advice_9 == memory_0[79: 16] && In_timestamp == memory_0[207: 144] && 4'd0 == memory_0[11: 8] && 1'b1 == memory_0[0: 0] && 6'b000000 == memory_0[7: 2] && 1'b0 == memory_0[1: 1];
wire [1:0] v1ba = 2'b00;
wire v1bb = v1ba == v123;
wire v1bc = v72 & v72 & v72 & v72;
wire v1bd = v121 & v1bb & v115 & v1bc;
wire v1be = Advice_12 == Advice_11;
wire v1bf = v14e == Advice_3;
wire v1c0 = v146 & v1b6 & v11f & v1b8 & v11 & v13 & v1b9 & v1bd & v7a & v78 & v127 & v14b & v14c & v1be & v14d & va2 & v1bf;
wire rnx2x15 = rnx2x14 || v1c0;
wire onx2x15 = onx2x14 || ( rnx2x14 && v1c0);
wire [31:0] v1c1 = v1b4 + v11c;
wire v1c2 = v1c1 == Advice_9;
wire [1:0] v1c3 = 2'b10;
wire v1c4 = v1c3 == v123;
wire v1c5 = Advice_7 == v13f;
wire v1c6 = v1c5;
wire v1c7 = v1c6 ^ v72;
wire v1c8 = Advice_12 == v13f;
wire v1c9 = v1c8;
wire v1ca = v1c9 ^ v72;
wire v1cb = v72 & v1c7 & v72 & v1ca;
wire v1cc = v121 & v1c4 & ved & v1cb;
wire v1cd = v154 & v14b & v1c2 & v13 & v11 & v1b9 & v1b8 & v1cc & v127 & v158 & v78 & v7a & v14c & v1be & v14d & va2 & v1bf;
wire rnx2x16 = rnx2x15 || v1cd;
wire onx2x16 = onx2x15 || ( rnx2x15 && v1cd);
wire [7:0] v1ce = instruction_bits[55: 48];
wire [7:0] pad_463 = (v1ce[7:7] == 1'b1) ?24'b111111111111111111111111 : 24'b000000000000000000000000;
wire [31:0] v1cf = { pad_463, v1ce };
wire v1d1 = v1cf == Advice_6;
wire [1:0] v1d2 = 2'b01;
wire v1d3 = v1d2 == v123;
wire v1d4 = v72 & v72 & v72 & v1ca;
wire v1d5 = v121 & v1d3 & vb3 & v1d4;
wire [31:0] v1d6 = v1b4 + v85;
wire v1d7 = v1d6 == Advice_9;
wire v1d8 = v1a4 & v127 & v1d1 & v1b9 & v1b8 & v14b & v11 & v13 & v1d5 & v7a & v78 & v1d7 & v14c & v1be & v14d & va2 & v1bf;
wire rnx2x17 = rnx2x16 || v1d8;
wire onx2x17 = onx2x16 || ( rnx2x16 && v1d8);
wire v1d9 = v87 == Advice_9;
wire [10:0] v1da = 11'b11010110101;
wire [10:0] v1db = instruction_bits[10: 0];
wire v1dc = v1da == v1db;
wire v1dd = v1dc & v1bb & vb3 & v1bc;
wire v1de = v13 & v1d1 & v78 & v1d9 & v1dd & v1b9 & v1a4 & v11 & v14b & v7a & v14d & va2 & v1bf;
wire rnx2x18 = rnx2x17 || v1de;
wire onx2x18 = onx2x17 || ( rnx2x17 && v1de);
wire [31:0] v1df = { 30'b000000000000000000000000000000, v15f };
wire [31:0] v1e1 = v17f << v1df;
wire [31:0] v1e2 = v1b3 + v1e1;
wire [31:0] v1e3 = v1e2 + v4;
wire v1e4 = v1e3 == Advice_9;
wire [10:0] v1e5 = 11'b11010110001;
wire v1e6 = v1e5 == v1db;
wire v1e8 = Advice_13 == v13f;
wire v1e9 = v1e8;
wire v1ea = v1e9 ^ v72;
wire v1eb = Advice_12 == v142;
wire v1ec = v1eb;
wire v1ed = v1ec ^ v72;
wire v1ee = v72 & v72 & v1ea & v1ed;
wire v1ef = v1e6 & v1bb & ved & v1ee;
wire v1f0 = v118 == Advice_12;
wire v1f1 = v15b == Advice_13;
wire v1f2 = Advice_13 == Advice_10;
wire v1f3 = v154 & v1e4 & v13 & v1ef & v1b9 & v158 & v1f0 & v1f1 & v78 & v7a & v159 & v11 & v14b & v14c & v1f2 & v1be & v14d & va2 & v1bf;
wire rnx2x19 = rnx2x18 || v1f3;
wire onx2x19 = onx2x18 || ( rnx2x18 && v1f3);
wire [7:0] v1f4 = instruction_bits[63: 56];
wire [7:0] pad_501 = (v1f4[7:7] == 1'b1) ?24'b111111111111111111111111 : 24'b000000000000000000000000;
wire [31:0] v1f5 = { pad_501, v1f4 };
wire v1f7 = v1f5 == Advice_6;
wire [31:0] v1f8 = v1e2 + va6;
wire v1f9 = v1f8 == Advice_9;
wire v1fa = Advice_7 == v12c;
wire v1fb = Advice_7 == v133;
wire v1fc = Advice_7 == v136;
wire v1fd = Advice_7 == v130;
wire v1fe = Advice_7 == v139;
wire v1ff = Advice_7 == v13c;
wire v200 = v1fa & v1fb & v1fc & v1fd & v1fe & v1ff;
wire v201 = v200 ^ v72;
wire v202 = v72 & v201 & v1ea & v72;
wire v203 = v1e6 & v1d3 & v71 & v202;
wire v204 = v1af & v1f7 & v1f9 & v203 & v1b9 & v14b & v1f1 & v1f0 & v13 & v159 & v11 & v78 & v7a & v14c & v1f2 & v1be & v14d & va2 & v1bf;
wire rnx2x20 = rnx2x19 || v204;
wire onx2x20 = onx2x19 || ( rnx2x19 && v204);
wire [31:0] v205 = v1e2 + v156;
wire v206 = v205 == Advice_9;
wire v207 = v1e6 & v1c4 & v16c & v202;
wire v208 = v172 & v176 & v206 & v11 & v1b9 & v13 & v1f0 & v1f1 & v159 & v7a & v78 & v14b & v207 & v14c & v1f2 & v1be & v14d & va2 & v1bf;
wire rnx2x21 = rnx2x20 || v208;
wire onx2x21 = onx2x20 || ( rnx2x20 && v208);
wire [31:0] v20a = ( Advice_14 == 2'd0) ? In_register_EDX :
	( Advice_14 == 2'd1) ? In_register_ESI :
	( Advice_14 == 2'd2) ? In_register_EBX : In_register_EDI;
wire [31:0] v20b = v20a << v1df;
wire [31:0] v20c = v6 + v20b;
wire [31:0] v20d = v20c + va6;
wire v20e = v20d == Advice_9;
wire v210 = instruction_bits[19: 19];
wire v20f = instruction_bits[21: 21];
wire [1:0] v211 = { v210 , v20f };
wire v213 = v211 == Advice_15;
wire [4:0] v214 = 5'b00101;
wire [4:0] v215 = instruction_bits[18: 14];
wire v216 = v214 == v215;
wire v217 = instruction_bits[20: 20];
wire v218 = v72 == v217;
wire v219 = v1e6 & v216 & v218 & v71 & v1bc;
wire v21a = Advice_15 == Advice_14;
wire v21b = v1f7 & v1af & v20e & v11 & v1b9 & v14b & v78 & v213 & v219 & v13 & v7a & v21a & v14d & va2 & v1bf;
wire rnx2x22 = rnx2x21 || v21b;
wire onx2x22 = onx2x21 || ( rnx2x21 && v21b);
wire [31:0] v21c = v1b4 + va6;
wire v21d = v21c == Advice_9;
wire [4:0] v21e = 5'b00111;
wire v21f = v21e == v111;
wire v220 = v1e6 & v1d3 & v21f & v71 & v1bc;
wire v221 = v1af & v1f0 & v21d & v220 & v13 & v11 & v159 & v14b & v1b9 & v7a & v78 & v1f7 & v14c & v1be & v14d & va2 & v1bf;
wire rnx2x23 = rnx2x22 || v221;
wire onx2x23 = onx2x22 || ( rnx2x22 && v221);
wire v222 = v72 & v72 & v72 & v1ed;
wire v223 = v1e6 & v1bb & v21f & ved & v222;
wire v224 = v154 & v1b6 & v13 & v11 & v158 & v1b9 & v1f0 & v14b & v223 & v7a & v78 & v159 & v14c & v1be & v14d & va2 & v1bf;
wire rnx2x24 = rnx2x23 || v224;
wire onx2x24 = onx2x23 || ( rnx2x23 && v224);
wire [31:0] v225 = v1b4 + v156;
wire v226 = v225 == Advice_9;
wire v227 = v1e6 & v1c4 & v21f & v16c & v1bc;
wire v228 = v226 & v14b & v11 & v13 & v176 & v159 & v172 & v1f0 & v227 & v7a & v78 & v1b9 & v14c & v1be & v14d & va2 & v1bf;
wire rnx2x25 = rnx2x24 || v228;
wire onx2x25 = onx2x24 || ( rnx2x24 && v228);
wire [31:0] v22a = ( Advice_16 == 3'd0) ? In_register_ESBASE :
	( Advice_16 == 3'd1) ? In_register_ESBASE :
	( Advice_16 == 3'd2) ? In_register_ESBASE :
	( Advice_16 == 3'd3) ? In_register_ESBASE :
	( Advice_16 == 3'd4) ? In_register_ESBASE :
	( Advice_16 == 3'd5) ? In_register_ESBASE :
	( Advice_16 == 3'd6) ? In_register_ESBASE : In_register_ESBASE;
wire [31:0] v22b = v22a + ve2;
wire [31:0] v22c = v22b + v7;
wire [31:0] v22d = v22c + va6;
wire v22e = v22d == Advice_9;
wire v22f = v1d2 == v15f;
wire v230 = v15e & v22f & v71 & v1cb;
wire v231 = Advice_12 == Advice_16;
wire v232 = v22e & v1f7 & v13 & v11 & v1f0 & v159 & v15c & v1b9 & v1af & v230 & v78 & v7a & v14c & v231 & v14d & va2 & v1bf;
wire rnx2x26 = rnx2x25 || v232;
wire onx2x26 = onx2x25 || ( rnx2x25 && v232);
wire [7:0] v233 = instruction_bits[47: 40];
wire [7:0] pad_564 = (v233[7:7] == 1'b1) ?24'b111111111111111111111111 : 24'b000000000000000000000000;
wire [31:0] v234 = { pad_564, v233 };
wire v236 = v234 == Advice_6;
wire v237 = instruction_bits[17: 17];
wire v238 = { v237 };
wire v23a = v238 == Advice_17;
wire [31:0] v23c = ( Advice_18 == 3'd0) ? In_register_EBX :
	( Advice_18 == 3'd1) ? In_register_EBX :
	( Advice_18 == 3'd2) ? In_register_EBP :
	( Advice_18 == 3'd3) ? In_register_EBP :
	( Advice_18 == 3'd4) ? In_register_ESI :
	( Advice_18 == 3'd5) ? In_register_EDI :
	( Advice_18 == 3'd6) ? In_register_EBP : In_register_EBX;
wire [31:0] v23d = v23c & ve3;
wire [31:0] v23e = v1b2 + v23d;
wire [31:0] v240 = ( Advice_19 == 1'd0) ? In_register_ESI : In_register_EDI;
wire [31:0] v241 = v240 & ve3;
wire [31:0] v242 = 32'b10000000000000000000000000000000;
wire [31:0] v244 = v241 << v242;
wire [31:0] v245 = v23e + v244;
wire [31:0] v246 = v245 + v17a;
wire [15:0] v247 = v246[15:0];
wire [31:0] v248 = { 16'b0000000000000000, v247 };
wire v249 = v248 == Advice_9;
wire v24b = v238 == Advice_20;
wire [15:0] v24c = 16'b1110011011010110;
wire v24d = v24c == v9b;
wire v24e = instruction_bits[18: 18];
wire v24f = vf == v24e;
wire v250 = Advice_20;
wire v251 = v250 ^ v72;
wire v252 = v72 & v251 & v72 & v72;
wire v253 = v24d & v24f & v22f & v9f & v252;
wire v254 = instruction_bits[16: 16];
wire v255 = { v254 };
wire v257 = v255 == Advice_21;
wire [2:0] v258 = { Advice_20 , v1ba };
wire v259 = v258 == Advice_18;
wire v25a = Advice_21 == Advice_19;
wire [2:0] v25b = { Advice_17 , v1ba };
wire v25c = v25b == Advice_11;
wire v25d = v19e & v236 & v13 & v23a & v7a & v78 & v249 & v1b9 & v24b & v11 & v15c & v253 & v257 & v259 & v25a & v25c & v14d & va2 & v1bf;
wire rnx2x27 = rnx2x26 || v25d;
wire onx2x27 = onx2x26 || ( rnx2x26 && v25d);
wire [7:0] v25e = instruction_bits[71: 64];
wire [7:0] pad_607 = (v25e[7:7] == 1'b1) ?24'b111111111111111111111111 : 24'b000000000000000000000000;
wire [31:0] v25f = { pad_607, v25e };
wire v261 = v25f == Advice_6;
wire [31:0] v262 = { 30'b000000000000000000000000000000, v168 };
wire [31:0] v264 = v17f << v262;
wire [31:0] v265 = v22b + v264;
wire [31:0] v266 = v265 + va;
wire v267 = v266 == Advice_9;
wire [18:0] v268 = 19'b0110010011010110001;
wire [18:0] v269 = instruction_bits[18: 0];
wire v26a = v268 == v269;
wire [47:0] v26b = 48'b000000000000000000000000000000000000000000000000;
wire [47:0] v26c = instruction_bits[119: 72];
wire v26d = v26b == v26c;
wire v26e = v72 & v72 & v1ea & v72;
wire v26f = v26a & v22f & v26d & v26e;
wire v270 = vde == Advice_12;
wire v271 = v164 == Advice_13;
wire [31:0] v272 = 32'b10010000000000000000000000000000;
wire [31:0] v273 = In_register_EIP + v272;
wire v274 = v273 == Out_register_EIP;
wire v275 = v12f & v132 & v135 & v138 & v13b & v13e & v141 & v144 & v274 & v42 & v45 & v48 & v4a & v4d & v50 & v53 & v97 & v5b & v98 & v60 & v63 & v66;
wire v276 = v12b & v275;
wire v277 = v261 & v267 & v11 & v26f & v270 & v15c & v13 & v177 & v1b9 & v271 & v276 & v78 & v7a & v14c & v1f2 & v231 & v14d & va2 & v1bf;
wire rnx2x28 = rnx2x27 || v277;
wire onx2x28 = onx2x27 || ( rnx2x27 && v277);
wire v278 = va8 == Advice_9;
wire [9:0] v279 = 10'b0010100111;
wire [9:0] v27a = instruction_bits[23: 14];
wire v27b = v279 == v27a;
wire v27c = v1e6 & v27b & v71 & v1bc;
wire v27d = v1f7 & v14b & v1af & v278 & v27c & v11 & v13 & v1b9 & v78 & v7a & v14d & va2 & v1bf;
wire rnx2x29 = rnx2x28 || v27d;
wire onx2x29 = onx2x28 || ( rnx2x28 && v27d);
wire [31:0] v27e = In_register_FSBASE + v4;
wire [31:0] v27f = v27e + v7;
wire [31:0] v280 = v27f + va6;
wire v281 = v280 == Advice_9;
wire [18:0] v282 = 19'b0010011011010110101;
wire v283 = v282 == v269;
wire v284 = v1ba == v15f;
wire v285 = v283 & v284 & v71 & v1bc;
wire v286 = v281 & v13 & v1b9 & v1af & v15c & v11 & v285 & v78 & v1f7 & v7a & v14d & va2 & v1bf;
wire rnx2x30 = rnx2x29 || v286;
wire onx2x30 = onx2x29 || ( rnx2x29 && v286);
wire [1:0] v287 = { v254 , v24e };
wire v289 = v287 == Advice_22;
wire [31:0] v28a = v22a + v20a;
wire [31:0] v28b = v28a + v7;
wire [31:0] v28c = v28b + v4;
wire v28d = v28c == Advice_9;
wire v28e = v72 == v237;
wire v28f = v15e & v28e & v284 & ved & v1bc;
wire v291 = v287 == Advice_23;
wire v292 = Advice_22 == Advice_14;
wire [2:0] v293 = { Advice_23 , vf };
wire v294 = v293 == Advice_16;
wire v295 = v154 & v158 & v11 & v1b9 & v13 & v289 & v15c & v28d & v28f & v7a & v78 & v291 & v292 & v294 & v14d & va2 & v1bf;
wire rnx2x31 = rnx2x30 || v295;
wire onx2x31 = onx2x30 || ( rnx2x30 && v295);
wire v296 = v1c3 == v15f;
wire v297 = v15e & v296 & v16c & v1cb;
wire [31:0] v298 = v22c + v156;
wire v299 = v298 == Advice_9;
wire v29a = v172 & v11 & v13 & v1b9 & v176 & v297 & v159 & v7a & v78 & v1f0 & v15c & v299 & v14c & v231 & v14d & va2 & v1bf;
wire rnx2x32 = rnx2x31 || v29a;
wire onx2x32 = onx2x31 || ( rnx2x31 && v29a);
wire [31:0] v29c = ( Advice_24 == 3'd0) ? In_register_FSBASE :
	( Advice_24 == 3'd1) ? In_register_FSBASE :
	( Advice_24 == 3'd2) ? In_register_FSBASE :
	( Advice_24 == 3'd3) ? In_register_FSBASE :
	( Advice_24 == 3'd4) ? In_register_FSBASE :
	( Advice_24 == 3'd5) ? In_register_FSBASE :
	( Advice_24 == 3'd6) ? In_register_FSBASE : In_register_FSBASE;
wire [31:0] v29d = v29c + ve2;
wire [31:0] v29e = v29d + v264;
wire [31:0] v29f = v29e + v174;
wire v2a0 = v29f == Advice_9;
wire [18:0] v2a1 = 19'b0010011011010110001;
wire v2a2 = v2a1 == v269;
wire v2a3 = v2a2 & v296 & v9f & v26e;
wire v2a4 = Advice_12 == Advice_24;
wire v2a5 = v19e & v236 & v271 & v11 & v7a & v78 & v1b9 & v270 & v13 & v15c & v2a0 & v177 & v2a3 & v14c & v1f2 & v2a4 & v14d & va2 & v1bf;
wire rnx2x33 = rnx2x32 || v2a5;
wire onx2x33 = onx2x32 || ( rnx2x32 && v2a5);
wire [31:0] v2a7 = ( Advice_25 == 2'd0) ? In_register_DSBASE :
	( Advice_25 == 2'd1) ? In_register_DSBASE :
	( Advice_25 == 2'd2) ? In_register_DSBASE : In_register_DSBASE;
wire [31:0] v2a9 = ( Advice_26 == 1'd0) ? In_register_EDI : In_register_EBX;
wire [31:0] v2aa = v2a9 & ve3;
wire [31:0] v2ab = v2a7 + v2aa;
wire [31:0] v2ac = v2ab + v7;
wire [31:0] v2ad = v2ac + v4;
wire [15:0] v2ae = v2ad[15:0];
wire [31:0] v2af = { 16'b0000000000000000, v2ae };
wire v2b0 = v2af == Advice_9;
wire [16:0] v2b1 = 17'b11100110110101101;
wire [16:0] v2b2 = instruction_bits[16: 0];
wire v2b3 = v2b1 == v2b2;
wire v2b4 = v72 == v24e;
wire v2b5 = v2b3 & v2b4 & v284 & ved & v1bc;
wire v2b6 = Advice_20 == Advice_26;
wire [1:0] v2b7 = { Advice_17 , vf };
wire v2b8 = v2b7 == Advice_25;
wire v2b9 = v2b0 & v154 & v13 & v158 & v1b9 & v11 & v15c & v2b5 & v7a & v78 & v24b & v23a & v2b6 & v2b8 & v14d & va2 & v1bf;
wire rnx2x34 = rnx2x33 || v2b9;
wire onx2x34 = onx2x33 || ( rnx2x33 && v2b9);
wire v2ba = v24d & v24f & v296 & v16c & v252;
wire [31:0] v2bb = v245 + v156;
wire [15:0] v2bc = v2bb[15:0];
wire [31:0] v2bd = { 16'b0000000000000000, v2bc };
wire v2be = v2bd == Advice_9;
wire v2bf = v176 & v172 & v2ba & v2be & v24b & v13 & v1b9 & v23a & v257 & v78 & v7a & v15c & v11 & v259 & v25a & v25c & v14d & va2 & v1bf;
wire rnx2x35 = rnx2x34 || v2bf;
wire onx2x35 = onx2x34 || ( rnx2x34 && v2bf);
wire [31:0] v2c0 = v245 + v4;
wire [15:0] v2c1 = v2c0[15:0];
wire [31:0] v2c2 = { 16'b0000000000000000, v2c1 };
wire v2c3 = v2c2 == Advice_9;
wire v2c4 = v24d & v24f & v284 & ved & v252;
wire v2c5 = v154 & v2c3 & v11 & v13 & v23a & v24b & v2c4 & v257 & v158 & v7a & v78 & v15c & v1b9 & v259 & v25a & v25c & v14d & va2 & v1bf;
wire rnx2x36 = rnx2x35 || v2c5;
wire onx2x36 = onx2x35 || ( rnx2x35 && v2c5);
wire [15:0] v2c6 = 16'b0000000111111111;
wire [15:0] v2c7 = vb8 + v2c6;
wire [15:0] v2c8 = 16'b0000000011111111;
wire v2c9 = v2c7 < v2c8;
wire v2ca = v2c9 == Out_register_CF;
wire v2cb = v2c9 == Out_register_OF;
wire v2cc = vc4 & v22 & v25 & vc5 & v31 & v34 & v37 & v3a & vac & v42 & v45 & v48 & v4a & v4d & v50 & v53 & v2ca & v5b & v2cb & v60 & v63 & v66;
wire v2cd = v1f8 == Advice_1;
wire [15:0] v2ce = 16'b0110111100110101;
wire v2cf = v2ce == v9b;
wire v2d0 = v72 & v1c7 & v72;
wire v2d1 = v2cf & vb3 & v2d0;
wire v2d2 = v118 == Advice_13;
wire v2d3 = v15b == Advice_7;
wire v2d4 = Advice_7 == Advice_10;
wire v2d5 = Advice_13 == Advice_11;
wire [7:0] pad_726 = (vd0[7:7] == 1'b1) ?8'b11111111 : 8'b00000000;
wire [15:0] v2d6 = { pad_726, vd0 };
wire [15:0] pad_727 = (v2d6[15:15] == 1'b1) ?48'b111111111111111111111111111111111111111111111111 : 48'b000000000000000000000000000000000000000000000000;
wire [63:0] v2d7 = { pad_727, v2d6 };
wire v2d8 = v2d7 == Advice_2;
wire [7:0] pad_729 = (vd4[7:7] == 1'b1) ?8'b11111111 : 8'b00000000;
wire [15:0] v2d9 = { pad_729, vd4 };
wire [15:0] pad_730 = (v2d9[15:15] == 1'b1) ?48'b111111111111111111111111111111111111111111111111 : 48'b000000000000000000000000000000000000000000000000;
wire [63:0] v2da = { pad_730, v2d9 };
wire v2db = v2da == Advice_3;
wire v2dc = v2cc & v2cd & v11 & v13 & vcf & v119 & v2d1 & v78 & v2d2 & v2d3 & v7a & vf0 & v2d4 & v2d5 & v2d8 & v2db;
wire rnx2x37 = rnx2x36 || v2dc;
wire onx2x37 = onx2x36 || ( rnx2x36 && v2dc);
wire [31:0] v2dd = ve2 << v262;
wire [31:0] v2de = v28a + v2dd;
wire [31:0] v2df = v2de + v4;
wire v2e0 = v2df == Advice_9;
wire v2e1 = instruction_bits[25: 25];
wire v2e2 = v72 == v2e1;
wire v2e3 = v26a & v284 & v2e2 & v16c & v26e;
wire v2e5 = instruction_bits[24: 24];
wire v2e4 = instruction_bits[26: 26];
wire [1:0] v2e6 = { v2e5 , v2e4 };
wire v2e7 = v2e6 == Advice_23;
wire v2e8 = v2e6 == Advice_22;
wire v2e9 = Advice_13 == Advice_5;
wire v2ea = v172 & v176 & v11 & v271 & v13 & v2e0 & v2e3 & v2e7 & v15c & v2e8 & v1b9 & v78 & v7a & v292 & v2e9 & v294 & v14d & va2 & v1bf;
wire rnx2x38 = rnx2x37 || v2ea;
wire onx2x38 = onx2x37 || ( rnx2x37 && v2ea);
wire v2eb = v12f & v132 & v135 & v138 & v13b & v13e & v141 & v144 & v274 & v42 & v45 & v48 & v4a & v4d & v50 & v53 & v58 & v5b & v5d & v60 & v63 & v66;
wire v2ec = v182 & v2eb;
wire [15:0] v2ed = instruction_bits[71: 56];
wire [15:0] pad_750 = (v2ed[15:15] == 1'b1) ?16'b1111111111111111 : 16'b0000000000000000;
wire [31:0] v2ee = { pad_750, v2ed };
wire v2f0 = v2ee == Advice_6;
wire v2f1 = v186 & v22f & v26d & v1cb;
wire v2f2 =  v69 == memory_0[15: 12] && Advice_9 == memory_0[79: 16] && In_timestamp == memory_0[207: 144] && 4'd0 == memory_0[11: 8] && 1'b1 == memory_0[0: 0] && 6'b000000 == memory_0[7: 2] && 1'b0 == memory_0[1: 1];
wire v2f3 = v7e == Advice_3;
wire v2f4 = v2ec & v1f0 & v2f0 & v7a & v2f1 & v78 & v15c & v13 & v159 & v21d & v11 & v2f2 & v14c & v1be & v14d & v188 & v18c & v2f3;
wire rnx2x39 = rnx2x38 || v2f4;
wire onx2x39 = onx2x38 || ( rnx2x38 && v2f4);
wire [31:0] v2f6 = ( Advice_27 == 3'd0) ? In_register_EAX :
	( Advice_27 == 3'd1) ? In_register_ECX :
	( Advice_27 == 3'd2) ? In_register_EDX :
	( Advice_27 == 3'd3) ? In_register_EBX :
	( Advice_27 == 3'd4) ? In_register_ESP :
	( Advice_27 == 3'd5) ? In_register_EBP :
	( Advice_27 == 3'd6) ? In_register_ESI : In_register_EDI;
wire [15:0] v2f7 = v2f6[31: 16];
wire [31:0] v2f8 = { v2f7 , v1b };
wire v2f9 = v2f8 == v12a;
wire [31:0] v2fa = 32'b01010000000000000000000000000000;
wire [31:0] v2fb = In_register_EIP + v2fa;
wire v2fc = v2fb == Out_register_EIP;
wire v2fd = v12f & v132 & v135 & v138 & v13b & v13e & v141 & v144 & v2fc & v42 & v45 & v48 & v4a & v4d & v50 & v53 & v58 & v5b & v5d & v60 & v63 & v66;
wire v2fe = v2f9 & v2fd;
wire [15:0] v2ff = instruction_bits[79: 64];
wire [15:0] pad_768 = (v2ff[15:15] == 1'b1) ?16'b1111111111111111 : 16'b0000000000000000;
wire [31:0] v300 = { pad_768, v2ff };
wire v302 = v300 == Advice_6;
wire [18:0] v303 = 19'b0110011010010110001;
wire v304 = v303 == v269;
wire [39:0] v305 = 40'b0000000000000000000000000000000000000000;
wire [39:0] v306 = instruction_bits[119: 80];
wire v307 = v305 == v306;
wire v308 = v304 & v22f & v307 & v26e;
wire [31:0] v309 = v1b3 + v264;
wire [31:0] v30a = v309 + va;
wire v30b = v30a == Advice_9;
wire v30c = Advice_4 == Advice_27;
wire v30d = v2fe & v302 & v13 & v2f2 & v177 & v11 & v15c & v270 & v271 & v78 & v7a & v308 & v30b & v14c & v1f2 & v1be & v14d & v30c & v18c & v2f3;
wire rnx2x40 = rnx2x39 || v30d;
wire onx2x40 = onx2x39 || ( rnx2x39 && v30d);
wire v30e = v186 & v28e & v284 & v16c & v1bc;
wire [31:0] v30f = v2a7 + v20a;
wire [31:0] v310 = v30f + v7;
wire [31:0] v311 = v310 + v4;
wire v312 = v311 == Advice_9;
wire [15:0] v313 = ve2[31: 16];
wire [31:0] v314 = { v313 , v1b };
wire v315 = v314 == v12a;
wire v316 = v315 & v183;
wire v317 = Advice_23 == Advice_25;
wire v318 = v13 & v17c & v30e & v312 & v15c & v11 & v289 & v316 & v2f2 & v291 & v78 & v7a & v292 & v317 & v14d & vf0 & v18c & v2f3;
wire rnx2x41 = rnx2x40 || v318;
wire onx2x41 = onx2x40 || ( rnx2x40 && v318);
wire v319 = v186 & v296 & v9f & v1d4;
wire v31a = v19a & v11 & v13 & v2f2 & v193 & v1f0 & v159 & v319 & v15c & v7a & v78 & v226 & v14c & v1be & v14d & v188 & v18c & v2f3;
wire rnx2x42 = rnx2x41 || v31a;
wire onx2x42 = onx2x41 || ( rnx2x41 && v31a);
wire v31b = v12f & v132 & v135 & v138 & v13b & v13e & v141 & v144 & vac & v42 & v45 & v48 & v4a & v4d & v50 & v53 & v58 & v5b & v5d & v60 & v63 & v66;
wire v31c = v2f9 & v31b;
wire [31:0] v31d = v309 + v174;
wire v31e = v31d == Advice_9;
wire [15:0] v31f = instruction_bits[55: 40];
wire [15:0] pad_800 = (v31f[15:15] == 1'b1) ?16'b1111111111111111 : 16'b0000000000000000;
wire [31:0] v320 = { pad_800, v31f };
wire v322 = v320 == Advice_6;
wire v323 = v304 & v296 & vb3 & v26e;
wire v324 = v31c & v31e & v11 & v322 & v15c & v2f2 & v270 & v13 & v271 & v78 & v7a & v177 & v323 & v14c & v1f2 & v1be & v14d & v30c & v18c & v2f3;
wire rnx2x43 = rnx2x42 || v324;
wire onx2x43 = onx2x42 || ( rnx2x42 && v324);
wire [4:0] v325 = 5'b00110;
wire v326 = v325 == ve9;
wire v327 = Advice_7 == v142;
wire v328 = v327;
wire v329 = v328 ^ v72;
wire v32a = v72 & v329 & v72 & v1ed;
wire v32b = v304 & v284 & v326 & v9f & v32a;
wire v32c = v193 & v1b6 & v2f2 & v270 & v15c & v32b & v7a & v13 & v78 & v19a & v11 & v177 & v14c & v1be & v14d & v188 & v18c & v2f3;
wire rnx2x44 = rnx2x43 || v32c;
wire onx2x44 = onx2x43 || ( rnx2x43 && v32c);
wire v32d = v12f & v132 & v135 & v138 & v13b & v13e & v141 & v144 & v2fc & v42 & v45 & v48 & v4a & v4d & v50 & v53 & v97 & v5b & v98 & v60 & v63 & v66;
wire v32e = v12b & v32d;
wire [31:0] v32f = instruction_bits[79: 48];
wire v331 = v32f == Advice_6;
wire v333 = instruction_bits[8: 8];
wire v332 = instruction_bits[10: 10];
wire [1:0] v334 = { v333 , v332 };
wire v335 = v334 == Advice_23;
wire [31:0] v336 = v310 + v85;
wire v337 = v336 == Advice_9;
wire v338 = v334 == Advice_22;
wire v339 = instruction_bits[9: 9];
wire v33a = v72 == v339;
wire v33b = v1a0 & v33a & v1d3 & v307 & v1bc;
wire v33c = v32e & v331 & v13 & v335 & v337 & v338 & v11 & v1b9 & v14b & v33b & v78 & v7a & v292 & v317 & v14d & va2 & v1bf;
wire rnx2x45 = rnx2x44 || v33c;
wire onx2x45 = onx2x44 || ( rnx2x44 && v33c);
wire v33d = v1a0 & v1bb & v9f & v1bc;
wire v33e = v14b & v19c & v19e & v11 & v1b6 & v1b9 & v127 & v33d & v1b8 & v7a & v78 & v13 & v14c & v1be & v14d & va2 & v1bf;
wire rnx2x46 = rnx2x45 || v33e;
wire onx2x46 = onx2x45 || ( rnx2x45 && v33e);
wire [10:0] v33f = 11'b10010110101;
wire v340 = v33f == v1db;
wire v341 = v340 & v1bb & v307 & v1bc;
wire v342 = v331 & v1d9 & v13 & v14b & v11 & v341 & v1b9 & v32e & v78 & v7a & v14d & va2 & v1bf;
wire rnx2x47 = rnx2x46 || v342;
wire onx2x47 = onx2x46 || ( rnx2x46 && v342);
wire v343 = v1a0 & v1c4 & vb3 & v1cb;
wire v344 = v1a4 & v11 & v1b9 & v13 & v343 & v1a5 & v127 & v14b & v1b8 & v7a & v78 & v1c2 & v14c & v1be & v14d & va2 & v1bf;
wire rnx2x48 = rnx2x47 || v344;
wire onx2x48 = onx2x47 || ( rnx2x47 && v344);
wire [10:0] v345 = 11'b10010110001;
wire v346 = v345 == v1db;
wire v347 = v346 & v1bb & vb3 & v1ee;
wire v348 = v1a4 & v1a5 & v1b9 & v1e4 & v11 & v13 & v1f0 & v7a & v78 & v159 & v14b & v347 & v1f1 & v14c & v1f2 & v1be & v14d & va2 & v1bf;
wire rnx2x49 = rnx2x48 || v348;
wire onx2x49 = onx2x48 || ( rnx2x48 && v348);
wire v349 = v346 & v1c4 & v71 & v26e;
wire v34a = v1af & v1aa & v11 & v1b9 & v7a & v78 & v349 & v206 & v1f1 & v1f0 & v13 & v159 & v14b & v14c & v1f2 & v1be & v14d & va2 & v1bf;
wire rnx2x50 = rnx2x49 || v34a;
wire onx2x50 = onx2x49 || ( rnx2x49 && v34a);
wire [31:0] v34b = 32'b11010000000000000000000000000000;
wire [31:0] v34c = In_register_EIP + v34b;
wire v34d = v34c == Out_register_EIP;
wire v34e = v12f & v132 & v135 & v138 & v13b & v13e & v141 & v144 & v34d & v42 & v45 & v48 & v4a & v4d & v50 & v53 & v97 & v5b & v98 & v60 & v63 & v66;
wire v34f = v12b & v34e;
wire [31:0] v350 = instruction_bits[87: 56];
wire v352 = v350 == Advice_6;
wire [31:0] v353 = instruction_bits[119: 88];
wire v354 = v4 == v353;
wire v355 = v346 & v1d3 & v354 & v26e;
wire v356 = v34f & v352 & v1f0 & v11 & v159 & v355 & v13 & v1f9 & v1f1 & v7a & v14b & v78 & v1b9 & v14c & v1f2 & v1be & v14d & va2 & v1bf;
wire rnx2x51 = rnx2x50 || v356;
wire onx2x51 = onx2x50 || ( rnx2x50 && v356);
wire v357 = v346 & v1d3 & v21f & v354 & v1bc;
wire v358 = v34f & v352 & v21d & v1b9 & v1f0 & v357 & v159 & v13 & v14b & v11 & v78 & v7a & v14c & v1be & v14d & va2 & v1bf;
wire rnx2x52 = rnx2x51 || v358;
wire onx2x52 = onx2x51 || ( rnx2x51 && v358);
wire v359 = v346 & v1bb & v21f & vb3 & v222;
wire v35a = v78 & v7a & v1b6 & v11 & v1b9 & v1f0 & v13 & v159 & v14b & v1a5 & v1a4 & v359 & v14c & v1be & v14d & va2 & v1bf;
wire rnx2x53 = rnx2x52 || v35a;
wire onx2x53 = onx2x52 || ( rnx2x52 && v35a);
wire v35b = v346 & v1c4 & v21f & v71 & v1bc;
wire v35c = v1af & v14b & v11 & v1aa & v226 & v159 & v13 & v1b9 & v1f0 & v7a & v78 & v35b & v14c & v1be & v14d & va2 & v1bf;
wire rnx2x54 = rnx2x53 || v35c;
wire onx2x54 = onx2x53 || ( rnx2x53 && v35c);
wire v35d = v346 & v216 & v354 & v26e;
wire [31:0] v35e = ve2 << v1df;
wire [31:0] v35f = v6 + v35e;
wire [31:0] v360 = v35f + va6;
wire v361 = v360 == Advice_9;
wire v362 = v11 & v13 & v1b9 & v352 & v7a & v1f1 & v14b & v34f & v35d & v361 & v78 & v2e9 & v14d & va2 & v1bf;
wire rnx2x55 = rnx2x54 || v362;
wire onx2x55 = onx2x54 || ( rnx2x54 && v362);
wire [31:0] v363 = instruction_bits[71: 40];
wire v365 = v363 == Advice_6;
wire [31:0] v367 = ( Advice_28 == 3'd0) ? In_register_DSBASE :
	( Advice_28 == 3'd1) ? In_register_DSBASE :
	( Advice_28 == 3'd2) ? In_register_SSBASE :
	( Advice_28 == 3'd3) ? In_register_SSBASE :
	( Advice_28 == 3'd4) ? In_register_DSBASE :
	( Advice_28 == 3'd5) ? In_register_DSBASE :
	( Advice_28 == 3'd6) ? In_register_SSBASE : In_register_DSBASE;
wire [31:0] v368 = v367 + v23d;
wire [31:0] v36a = ( Advice_29 == 3'd0) ? In_register_ESI :
	( Advice_29 == 3'd1) ? In_register_EDI :
	( Advice_29 == 3'd2) ? In_register_ESI :
	( Advice_29 == 3'd3) ? In_register_EDI :
	( Advice_29 == 3'd4) ? v4 :
	( Advice_29 == 3'd5) ? v4 :
	( Advice_29 == 3'd6) ? v4 : v4;
wire [31:0] v36b = v36a & ve3;
wire [31:0] v36c = v36b << v242;
wire [31:0] v36d = v368 + v36c;
wire [31:0] v36e = v36d + v17a;
wire [15:0] v36f = v36e[15:0];
wire [31:0] v370 = { 16'b0000000000000000, v36f };
wire v371 = v370 == Advice_9;
wire v372 = v1a7 & v22f & v26d & v1bc;
wire v373 = Advice_7 == Advice_18;
wire v374 = Advice_13 == Advice_29;
wire v375 = Advice_12 == Advice_28;
wire v376 = v365 & v13 & v1b9 & v11 & v1f0 & v2d2 & v276 & v159 & v371 & v15c & v7a & v78 & v372 & v373 & v374 & v375 & v14d & va2 & v1bf;
wire rnx2x56 = rnx2x55 || v376;
wire onx2x56 = onx2x55 || ( rnx2x55 && v376);
wire [15:0] v377 = 16'b0110010010010110;
wire v378 = v377 == v9b;
wire v379 = v378 & v22f & v354 & v1cb;
wire v37a = v34f & v22e & v11 & v13 & v1b9 & v15c & v352 & v379 & v7a & v78 & v159 & v1f0 & v14c & v231 & v14d & va2 & v1bf;
wire rnx2x57 = rnx2x56 || v37a;
wire onx2x57 = onx2x56 || ( rnx2x56 && v37a);
wire [31:0] v37b = v29d + v7;
wire [31:0] v37c = v37b + v4;
wire v37d = v37c == Advice_9;
wire [15:0] v37e = 16'b0010011010010110;
wire v37f = v37e == v9b;
wire v380 = v37f & v284 & vb3 & v1bc;
wire v381 = v1a4 & v1a5 & v11 & v1b9 & v1f0 & v159 & v37d & v13 & v15c & v78 & v7a & v380 & v14c & v2a4 & v14d & va2 & v1bf;
wire rnx2x58 = rnx2x57 || v381;
wire onx2x58 = onx2x57 || ( rnx2x57 && v381);
wire [31:0] v383 = ( Advice_30 == 3'd0) ? In_register_GSBASE :
	( Advice_30 == 3'd1) ? In_register_GSBASE :
	( Advice_30 == 3'd2) ? In_register_GSBASE :
	( Advice_30 == 3'd3) ? In_register_GSBASE :
	( Advice_30 == 3'd4) ? In_register_GSBASE :
	( Advice_30 == 3'd5) ? In_register_GSBASE :
	( Advice_30 == 3'd6) ? In_register_GSBASE : In_register_GSBASE;
wire [31:0] v384 = v383 + ve2;
wire [31:0] v385 = v20a << v262;
wire [31:0] v386 = v384 + v385;
wire [31:0] v387 = v386 + v174;
wire v388 = v387 == Advice_9;
wire [18:0] v389 = 19'b1010011010010110001;
wire v38a = v389 == v269;
wire v38b = instruction_bits[28: 28];
wire v38c = v72 == v38b;
wire v38d = v38a & v296 & v38c & v26d & v1bc;
wire v38f = instruction_bits[27: 27];
wire v38e = instruction_bits[29: 29];
wire [1:0] v390 = { v38f , v38e };
wire v391 = v390 == Advice_15;
wire v392 = Advice_12 == Advice_30;
wire v393 = v276 & v15c & v388 & v11 & v13 & v365 & v1b9 & v38d & v270 & v78 & v7a & v391 & v177 & v14c & v21a & v392 & v14d & va2 & v1bf;
wire rnx2x59 = rnx2x58 || v393;
wire onx2x59 = onx2x58 || ( rnx2x58 && v393);
wire [9:0] v394 = 10'b0010100101;
wire v395 = v394 == v27a;
wire v396 = v346 & v395 & v354 & v1bc;
wire v397 = v34f & v352 & v278 & v11 & v13 & v78 & v1b9 & v14b & v396 & v7a & v14d & va2 & v1bf;
wire rnx2x60 = rnx2x59 || v397;
wire onx2x60 = onx2x59 || ( rnx2x59 && v397);
wire [31:0] v398 = v29c + v20a;
wire [31:0] v399 = v398 + v7;
wire [31:0] v39a = v399 + v156;
wire v39b = v39a == Advice_9;
wire v39c = v37f & v28e & v296 & v71 & v1bc;
wire v39d = v293 == Advice_24;
wire v39e = v1af & v1b9 & v11 & v1aa & v39b & v39c & v291 & v13 & v289 & v15c & v78 & v7a & v292 & v39d & v14d & va2 & v1bf;
wire rnx2x61 = rnx2x60 || v39e;
wire onx2x61 = onx2x60 || ( rnx2x60 && v39e);
wire [16:0] v39f = 17'b11100110100101101;
wire v3a0 = v39f == v2b2;
wire v3a1 = v3a0 & v2b4 & v284 & vb3 & v1bc;
wire v3a2 = v15c & v1a5 & v11 & v13 & v1a4 & v1b9 & v24b & v2b0 & v23a & v3a1 & v78 & v7a & v2b6 & v2b8 & v14d & va2 & v1bf;
wire rnx2x62 = rnx2x61 || v3a2;
wire onx2x62 = onx2x61 || ( rnx2x61 && v3a2);
wire v3a3 = v1a7 & v296 & v71 & v1bc;
wire [31:0] v3a4 = v36d + v156;
wire [15:0] v3a5 = v3a4[15:0];
wire [31:0] v3a6 = { 16'b0000000000000000, v3a5 };
wire v3a7 = v3a6 == Advice_9;
wire v3a8 = v1aa & v3a3 & v1b9 & v1f0 & v1af & v11 & v15c & v13 & v2d2 & v7a & v78 & v159 & v3a7 & v373 & v374 & v375 & v14d & va2 & v1bf;
wire rnx2x63 = rnx2x62 || v3a8;
wire onx2x63 = onx2x62 || ( rnx2x62 && v3a8);
wire [31:0] v3a9 = 32'b00110000000000000000000000000000;
wire [31:0] v3aa = In_register_EIP + v3a9;
wire v3ab = v3aa == Out_register_EIP;
wire v3ac = v12f & v132 & v135 & v138 & v13b & v13e & v141 & v144 & v3ab & v42 & v45 & v48 & v4a & v4d & v50 & v53 & v97 & v5b & v98 & v60 & v63 & v66;
wire v3ad = v12b & v3ac;
wire [31:0] v3ae = instruction_bits[95: 64];
wire v3b0 = v3ae == Advice_6;
wire [18:0] v3b1 = 19'b0110110010010110001;
wire v3b2 = v3b1 == v269;
wire [23:0] v3b3 = 24'b000000000000000000000000;
wire [23:0] v3b4 = instruction_bits[119: 96];
wire v3b5 = v3b3 == v3b4;
wire v3b6 = v3b2 & v22f & v3b5 & v26e;
wire [31:0] v3b8 = ( Advice_31 == 3'd0) ? In_register_SSBASE :
	( Advice_31 == 3'd1) ? In_register_SSBASE :
	( Advice_31 == 3'd2) ? In_register_SSBASE :
	( Advice_31 == 3'd3) ? In_register_SSBASE :
	( Advice_31 == 3'd4) ? In_register_SSBASE :
	( Advice_31 == 3'd5) ? In_register_SSBASE :
	( Advice_31 == 3'd6) ? In_register_SSBASE : In_register_SSBASE;
wire [31:0] v3b9 = v3b8 + ve2;
wire [31:0] v3ba = v3b9 + v264;
wire [31:0] v3bb = v3ba + va;
wire v3bc = v3bb == Advice_9;
wire v3bd = Advice_12 == Advice_31;
wire v3be = v3ad & v3b0 & v13 & v3b6 & v11 & v270 & v177 & v271 & v15c & v3bc & v1b9 & v78 & v7a & v14c & v1f2 & v3bd & v14d & va2 & v1bf;
wire rnx2x64 = rnx2x63 || v3be;
wire onx2x64 = onx2x63 || ( rnx2x63 && v3be);
wire [31:0] v3bf = In_register_GSBASE + v4;
wire [31:0] v3c0 = v3bf + v7;
wire [31:0] v3c1 = v3c0 + va6;
wire v3c2 = v3c1 == Advice_9;
wire [18:0] v3c3 = 19'b1010011010010110101;
wire v3c4 = v3c3 == v269;
wire v3c5 = v3c4 & v284 & v354 & v1bc;
wire v3c6 = v34f & v352 & v3c2 & v15c & v1b9 & v78 & v11 & v3c5 & v13 & v7a & v14d & va2 & v1bf;
wire rnx2x65 = rnx2x64 || v3c6;
wire onx2x65 = onx2x64 || ( rnx2x64 && v3c6);
wire v3c7 = v255 == Advice_17;
wire [31:0] v3c8 = v2a7 + v241;
wire [31:0] v3c9 = v3c8 + v7;
wire [31:0] v3ca = v3c9 + v4;
wire [15:0] v3cb = v3ca[15:0];
wire [31:0] v3cc = { 16'b0000000000000000, v3cb };
wire v3cd = v3cc == Advice_9;
wire v3ce = v255 == Advice_20;
wire [1:0] v3cf = instruction_bits[18: 17];
wire v3d0 = v1d2 == v3cf;
wire v3d1 = v1a7 & v3d0 & v284 & vb3 & v1bc;
wire v3d2 = Advice_20 == Advice_19;
wire v3d3 = v1a4 & v11 & v13 & v78 & v7a & v1a5 & v1b9 & v3c7 & v15c & v3cd & v3ce & v3d1 & v3d2 & v2b8 & v14d & va2 & v1bf;
wire rnx2x66 = rnx2x65 || v3d3;
wire onx2x66 = onx2x65 || ( rnx2x65 && v3d3);
wire [31:0] v3d5 = 32'b00000000000000000000000000000000;
wire [31:0] v3d6 = ( Advice_32 == 1'd0) ? v3d5 : In_register_EBP;
wire [31:0] v3d7 = v3d6 & ve3;
wire [31:0] v3d8 = v1b2 + v3d7;
wire [31:0] v3d9 = v3d8 + v244;
wire [31:0] v3da = v3d9 + v4;
wire [15:0] v3db = v3da[15:0];
wire [31:0] v3dc = { 16'b0000000000000000, v3db };
wire v3dd = v3dc == Advice_9;
wire v3de = Advice_32 == vf;
wire v3df = v3de;
wire v3e0 = v3df ^ v72;
wire v3e1 = v72 & v3e0 & v72 & v72;
wire v3e2 = v1a7 & v24f & v284 & vb3 & v3e1;
wire v3e3 = Advice_20 == Advice_32;
wire v3e4 = v1a4 & v1a5 & v11 & v13 & v15c & v1b9 & v23a & v3dd & v3e2 & v7a & v78 & v24b & v257 & v3e3 & v25a & v25c & v14d & va2 & v1bf;
wire rnx2x67 = rnx2x66 || v3e4;
wire onx2x67 = onx2x66 || ( rnx2x66 && v3e4);
wire [31:0] v3e5 = v384 + v264;
wire [31:0] v3e6 = v3e5 + v4;
wire v3e7 = v3e6 == Advice_9;
wire v3e8 = v72 & v329 & v1ea & v1ed;
wire v3e9 = v38a & v284 & v71 & v3e8;
wire v3ea = v1af & v3e7 & v11 & v13 & v1b9 & v3e9 & v271 & v15c & v1aa & v7a & v78 & v270 & v177 & v14c & v1f2 & v392 & v14d & va2 & v1bf;
wire rnx2x68 = rnx2x67 || v3ea;
wire onx2x68 = onx2x67 || ( rnx2x67 && v3ea);
wire v3eb = vc4 & v22 & v25 & vc5 & v31 & v34 & v37 & v3a & v10d & v42 & v45 & v48 & v4a & v4d & v50 & v53 & v2ca & v5b & v2cb & v60 & v63 & v66;
wire [31:0] v3ec = v30f + v35e;
wire [31:0] v3ed = v3ec + v4;
wire v3ee = v3ed == Advice_1;
wire v3ef = v287 == Advice_15;
wire v3f1 = v287 == Advice_33;
wire [15:0] v3f2 = 16'b0110111100110100;
wire v3f3 = v3f2 == v9b;
wire v3f4 = v3f3 & v28e & v115 & v2d0;
wire v3f5 = Advice_33 == Advice_14;
wire v3f6 = Advice_15 == Advice_25;
wire v3f7 = v3eb & v3ee & v11 & vcf & v3ef & v2d3 & v13 & v3f1 & v3f4 & v78 & v7a & v3f5 & v14c & v3f6 & v2d8 & v2db;
wire rnx2x69 = rnx2x68 || v3f7;
wire onx2x69 = onx2x68 || ( rnx2x68 && v3f7);
wire v3f8 = v22d == Advice_1;
wire [15:0] v3f9 = 16'b0110010001101111;
wire v3fa = v3f9 == v9b;
wire [4:0] v3fb = 5'b10101;
wire v3fc = v3fb == v111;
wire v3fd = v140;
wire v3fe = v3fd ^ v72;
wire v3ff = v3fe & v72 & v1ea;
wire v400 = v3fa & v3fc & vb3 & v3ff;
wire v401 = Advice_13 == Advice_16;
wire v402 = v3f8 & v13 & vcf & v11 & v119 & v7a & v2d2 & v78 & v2cc & v400 & vf0 & v401 & v2d8 & v2db;
wire rnx2x70 = rnx2x69 || v402;
wire onx2x70 = onx2x69 || ( rnx2x69 && v402);
wire v403 = v360 == Advice_1;
wire [18:0] v404 = 19'b0110111100110100101;
wire v405 = v404 == v269;
wire v406 = v405 & vb3 & v2d0;
wire v407 = v11 & vcf & v13 & v2d3 & v403 & v406 & v2cc & v78 & v7a & v14c & v2d8 & v2db;
wire rnx2x71 = rnx2x70 || v407;
wire onx2x71 = onx2x70 || ( rnx2x70 && v407);
wire v408 = v3dc == Advice_1;
wire [15:0] v409 = 16'b1110011001101111;
wire v40a = v409 == v9b;
wire [5:0] v40b = 6'b010100;
wire [5:0] v40c = instruction_bits[23: 18];
wire v40d = v40b == v40c;
wire v40e = v3e0 & v72 & v72;
wire v40f = v40a & v40d & v115 & v40e;
wire v410 = v238 == Advice_21;
wire v412 = v238 == Advice_34;
wire v413 = Advice_34 == Advice_32;
wire [2:0] v414 = { Advice_21 , v1ba };
wire v415 = v414 == Advice_11;
wire v416 = v3eb & v11 & v13 & vcf & v408 & v7a & v40f & v410 & v3ce & v412 & v78 & v413 & v3d2 & v415 & v2d8 & v2db;
wire rnx2x72 = rnx2x71 || v416;
wire onx2x72 = onx2x71 || ( rnx2x71 && v416);
wire [31:0] v417 = v3d9 + v156;
wire [15:0] v418 = v417[15:0];
wire [31:0] v419 = { 16'b0000000000000000, v418 };
wire v41a = v419 == Advice_1;
wire v41b = vc4 & v22 & v25 & vc5 & v31 & v34 & v37 & v3a & vdb & v42 & v45 & v48 & v4a & v4d & v50 & v53 & v2ca & v5b & v2cb & v60 & v63 & v66;
wire [5:0] v41c = 6'b010110;
wire v41d = v41c == v40c;
wire v41e = v40a & v41d & ved & v40e;
wire v41f = v41a & v11 & v13 & v412 & v41b & v410 & v7a & v41e & vcf & v3ce & v78 & v413 & v3d2 & v415 & v2d8 & v2db;
wire rnx2x73 = rnx2x72 || v41f;
wire onx2x73 = onx2x72 || ( rnx2x72 && v41f);
wire [31:0] v420 = v30f + v2dd;
wire [31:0] v421 = v420 + v4;
wire v422 = v421 == Advice_1;
wire v423 = v2e6 == Advice_15;
wire v424 = v2e6 == Advice_33;
wire [23:0] v425 = 24'b011001101110111100110100;
wire v426 = v425 == vaf;
wire v427 = v426 & v2e2 & ved & v2d0;
wire v428 = v164 == Advice_7;
wire v429 = vdc & v13 & v422 & v423 & v11 & v424 & v427 & v78 & v428 & v6b & v7a & v3f5 & v14c & v3f6 & v7f & v83;
wire rnx2x74 = rnx2x73 || v429;
wire onx2x74 = onx2x73 || ( rnx2x73 && v429);
wire v42a = vfc == Advice_13;
wire v42b = v1d6 == Advice_1;
wire v42c = v3fb == v101;
wire v42d = v100 & v42c & v9f & v3ff;
wire v42e = v99 & v13 & v8a & v42a & vfd & v42b & v11 & v42d & v78 & v7a & vf0 & v2d5 & va2 & va4;
wire rnx2x75 = rnx2x74 || v42e;
wire onx2x75 = onx2x74 || ( rnx2x74 && v42e);
wire v42f = v1b5 == Advice_1;
wire [4:0] v430 = 5'b10100;
wire v431 = v430 == v101;
wire v432 = v100 & v431 & v105 & v73;
wire v433 = vf9 & v42f & v8a & vfd & v42a & v11 & v13 & v7a & v432 & v78 & vf0 & v2d5 & va2 & va4;
wire rnx2x76 = rnx2x75 || v433;
wire onx2x76 = onx2x75 || ( rnx2x75 && v433);
wire [31:0] v434 = v310 + v11c;
wire v435 = v434 == Advice_1;
wire v436 = v334 == Advice_15;
wire [4:0] v437 = 5'b10110;
wire v438 = v437 == v101;
wire v439 = v100 & v33a & v438 & v115 & v73;
wire v43a = v334 == Advice_33;
wire v43b = v10e & v13 & v435 & v11 & v8a & v436 & v7a & v439 & v43a & v78 & v3f5 & v3f6 & va2 & va4;
wire rnx2x77 = rnx2x76 || v43b;
wire onx2x77 = onx2x76 || ( rnx2x76 && v43b);
wire v43c = v211 == Advice_22;
wire [31:0] v43d = v1b3 + v20b;
wire [31:0] v43e = v43d + v156;
wire v43f = v43e == Advice_1;
wire [15:0] v440 = 16'b1110111100110110;
wire v441 = v440 == v9b;
wire v442 = v12d & v134 & v137 & v131 & v13a & v13d;
wire v443 = v442 ^ v72;
wire v444 = v443 & v72 & v72;
wire v445 = v441 & v218 & ved & v444;
wire v446 = v8b & v22 & v25 & v8f & v31 & v34 & v37 & v3a & vdb & v42 & v45 & v48 & v4a & v4d & v50 & v53 & v97 & v5b & v98 & v60 & v63 & v66;
wire v447 = v11 & v119 & v78 & v43c & v43f & v13 & v2d2 & v445 & v446 & v8a & v7a & vf0 & v292 & v2d5 & va2 & va4;
wire rnx2x78 = rnx2x77 || v447;
wire onx2x78 = onx2x77 || ( rnx2x77 && v447);
wire [15:0] v448 = 16'b1110111100110100;
wire v449 = v448 == v9b;
wire v44a = v449 & v28e & v21f & v115 & v73;
wire v44b = v311 == Advice_1;
wire v44c = v13 & v11 & v8a & v3ef & v10e & v44a & v78 & v3f1 & v44b & v7a & v3f5 & v3f6 & va2 & va4;
wire rnx2x79 = rnx2x78 || v44c;
wire onx2x79 = onx2x78 || ( rnx2x78 && v44c);
wire v44d = v225 == Advice_1;
wire v44e = v441 & v21f & ved & v73;
wire v44f = v446 & v11 & v44d & v13 & v8a & v119 & v78 & v7a & v2d2 & v44e & vf0 & v2d5 & va2 & va4;
wire rnx2x80 = rnx2x79 || v44f;
wire onx2x80 = onx2x79 || ( rnx2x79 && v44f);
wire v450 = v8b & v22 & v25 & v8f & v31 & v34 & v37 & v3a & v3f & v42 & v45 & v48 & v4a & v4d & v50 & v53 & v97 & v5b & v98 & v60 & v63 & v66;
wire [31:0] v451 = v29e + va;
wire v452 = v451 == Advice_1;
wire v453 = vde == Advice_13;
wire [23:0] v454 = 24'b001001101110111100110101;
wire v455 = v454 == vaf;
wire v456 = v455 & v71 & v2d0;
wire v457 = Advice_13 == Advice_24;
wire v458 = v450 & v452 & v13 & v8a & v11 & v428 & v453 & v78 & ve0 & v456 & v7a & vf0 & v2d4 & v457 & va2 & va4;
wire rnx2x81 = rnx2x80 || v458;
wire onx2x81 = onx2x80 || ( rnx2x80 && v458);
wire v459 = v8b & v22 & v25 & v8f & v31 & v34 & v37 & v3a & v170 & v42 & v45 & v48 & v4a & v4d & v50 & v53 & v97 & v5b & v98 & v60 & v63 & v66;
wire v45a = v248 == Advice_1;
wire [5:0] v45b = 6'b010101;
wire v45c = v45b == v40c;
wire v45d = Advice_34;
wire v45e = v45d ^ v72;
wire v45f = v45e & v72 & v72;
wire v460 = v110 & v45c & v16c & v45f;
wire [2:0] v461 = { Advice_34 , v1ba };
wire v462 = v461 == Advice_18;
wire v463 = v11 & v13 & v8a & v459 & v45a & v410 & v3ce & v460 & v78 & v412 & v7a & v462 & v3d2 & v415 & va2 & va4;
wire rnx2x82 = rnx2x81 || v463;
wire onx2x82 = onx2x81 || ( rnx2x81 && v463);
wire [31:0] v464 = v3ba + v174;
wire v465 = v464 == Advice_1;
wire [23:0] v466 = 24'b011011001110111100110110;
wire v467 = v466 == vaf;
wire v468 = v467 & v16c & v2d0;
wire v469 = Advice_13 == Advice_31;
wire v46a = v465 & v11 & v459 & v13 & v8a & v453 & v428 & ve0 & v468 & v78 & v7a & vf0 & v2d4 & v469 & va2 & va4;
wire rnx2x83 = rnx2x82 || v46a;
wire onx2x83 = onx2x82 || ( rnx2x82 && v46a);
wire v46b = v2af == Advice_1;
wire [16:0] v46c = 17'b11100110111011111;
wire v46d = v46c == v2b2;
wire [5:0] v46e = 6'b110100;
wire v46f = v46e == v40c;
wire v470 = v46d & v46f & v115 & v73;
wire v471 = Advice_34 == Advice_26;
wire [1:0] v472 = { Advice_21 , vf };
wire v473 = v472 == Advice_25;
wire v474 = v46b & v11 & v10e & v8a & v13 & v470 & v412 & v78 & v410 & v7a & v471 & v473 & va2 & va4;
wire rnx2x84 = rnx2x83 || v474;
wire onx2x84 = onx2x83 || ( rnx2x83 && v474);
wire [63:0] v475 = 64'b1111111111111111111111111111111100000000000000000000000000000000;
wire v476 = v19 > v475;
wire v477 = v476 == Out_register_CF;
wire v478 = v476 == Out_register_OF;
wire v479 = v8b & v22 & v25 & v8f & v31 & v34 & v37 & v3a & vf8 & v42 & v45 & v48 & v4a & v4d & v50 & v53 & v477 & v5b & v478 & v60 & v63 & v66;
wire v47a = v21e == v101;
wire v47b = v100 & v47a & v105 & vee;
wire [63:0] v47c = { 32'b00000000000000000000000000000000, In_register_EAX };
wire v47d = v47c == Advice_2;
wire [63:0] v47e = { 32'b00000000000000000000000000000000, Advice_1 };
wire v47f = v47e == Advice_3;
wire v480 = vfa & vfd & v479 & v78 & v11 & v13 & v47b & v7a & vf0 & v47d & v47f;
wire rnx2x85 = rnx2x84 || v480;
wire onx2x85 = onx2x84 || ( rnx2x84 && v480);
wire [15:0] v481 = 16'b0110110011101111;
wire v482 = v481 == v9b;
wire v483 = v482 & v21f & v115 & vee;
wire v484 = v8b & v22 & v25 & v8f & v31 & v34 & v37 & v3a & v10d & v42 & v45 & v48 & v4a & v4d & v50 & v53 & v477 & v5b & v478 & v60 & v63 & v66;
wire v485 = vfa & v11 & v483 & v13 & v78 & v484 & v119 & v7a & vf0 & v47d & v47f;
wire rnx2x86 = rnx2x85 || v485;
wire onx2x86 = onx2x85 || ( rnx2x85 && v485);
wire [7:0] v486 = 8'b01101111;
wire v487 = v486 == vff;
wire v488 = v214 == v101;
wire v489 = v72 & v72 & v1ea;
wire v48a = v487 & v488 & v9f & v489;
wire v48b = v42b & vca & v11 & v13 & vcf & v48a & v7a & v42a & vfd & v78 & vf0 & v2d5 & vd3 & vd7;
wire rnx2x87 = rnx2x86 || v48b;
wire onx2x87 = onx2x86 || ( rnx2x86 && v48b);
wire [31:0] v48c = v43d + v4;
wire v48d = v48c == Advice_1;
wire v48e = vc4 & v22 & v25 & vc5 & v31 & v34 & v37 & v3a & v10d & v42 & v45 & v48 & v4a & v4d & v50 & v53 & vc8 & v5b & vc9 & v60 & v63 & v66;
wire [15:0] v48f = 16'b0110111100100100;
wire v490 = v48f == v9b;
wire v491 = Advice_13 == v142;
wire v492 = v491;
wire v493 = v492 ^ v72;
wire v494 = v72 & v72 & v493;
wire v495 = v490 & v218 & v115 & v494;
wire v496 = v48d & v11 & v13 & vcf & v2d2 & v43c & v48e & v119 & v78 & v495 & v7a & vf0 & v292 & v2d5 & vd3 & vd7;
wire rnx2x88 = rnx2x87 || v496;
wire onx2x88 = onx2x87 || ( rnx2x87 && v496);
wire v497 = vc4 & v22 & v25 & vc5 & v31 & v34 & v37 & v3a & vac & v42 & v45 & v48 & v4a & v4d & v50 & v53 & vc8 & v5b & vc9 & v60 & v63 & v66;
wire [31:0] v498 = v43d + va6;
wire v499 = v498 == Advice_1;
wire [15:0] v49a = 16'b0110111100100101;
wire v49b = v49a == v9b;
wire v49c = v49b & v218 & vb3 & v73;
wire v49d = v497 & v13 & v2d2 & vcf & v43c & v499 & v11 & v49c & v119 & v78 & v7a & vf0 & v292 & v2d5 & vd3 & vd7;
wire rnx2x89 = rnx2x88 || v49d;
wire onx2x89 = onx2x88 || ( rnx2x88 && v49d);
wire v49e = v21c == Advice_1;
wire [15:0] v49f = 16'b0110011001101111;
wire v4a0 = v49f == v9b;
wire v4a1 = v214 == v111;
wire v4a2 = v4a0 & v4a1 & vb3 & v3ff;
wire v4a3 = v11 & v49e & v13 & v497 & vcf & v7a & v2d2 & v78 & v119 & v4a2 & vf0 & v2d5 & vd3 & vd7;
wire rnx2x90 = rnx2x89 || v4a3;
wire onx2x90 = onx2x89 || ( rnx2x89 && v4a3);
wire [18:0] v4a4 = 19'b0110111100100100101;
wire v4a5 = v4a4 == v269;
wire v4a6 = v4a5 & vb3 & v2d0;
wire v4a7 = v11 & v13 & vcf & v2d3 & v4a6 & v497 & v78 & v403 & v7a & v14c & vd3 & vd7;
wire rnx2x91 = rnx2x90 || v4a7;
wire onx2x91 = onx2x90 || ( rnx2x90 && v4a7);
wire v4a8 = vc4 & v22 & v25 & vc5 & v31 & v34 & v37 & v3a & vdb & v42 & v45 & v48 & v4a & v4d & v50 & v53 & vc8 & v5b & vc9 & v60 & v63 & v66;
wire [23:0] v4a9 = 24'b011001100110111100100100;
wire v4aa = v4a9 == vaf;
wire v4ab = v4aa & v2e2 & ved & v2d0;
wire v4ac = v4a8 & v13 & vcf & v428 & v422 & v11 & v4ab & v78 & v423 & v424 & v7a & v3f5 & v14c & v3f6 & vd3 & vd7;
wire rnx2x92 = rnx2x91 || v4ac;
wire onx2x92 = onx2x91 || ( rnx2x91 && v4ac);
wire v4ad = v325 == v101;
wire v4ae = v100 & v33a & v4ad & v115 & v73;
wire [63:0] v4af = { 32'b00000000000000000000000000000000, v7b };
wire v4b0 = v4af == Advice_2;
wire v4b1 = v47c == Advice_3;
wire v4b2 = v484 & v7a & v43a & v13 & v4ae & v435 & v11 & v78 & v8a & v436 & v3f5 & v3f6 & v4b0 & v4b1;
wire rnx2x93 = rnx2x92 || v4b2;
wire onx2x93 = onx2x92 || ( rnx2x92 && v4b2);
wire [4:0] v4b3 = 5'b00100;
wire v4b4 = v4b3 == v101;
wire v4b5 = v100 & v4b4 & v105 & v73;
wire v4b6 = v42f & v11 & v13 & v8a & v42a & v4b5 & vfd & v78 & v479 & v7a & vf0 & v2d5 & v4b0 & v4b1;
wire rnx2x94 = rnx2x93 || v4b6;
wire onx2x94 = onx2x93 || ( rnx2x93 && v4b6);
wire v4b7 = v205 == Advice_1;
wire [15:0] v4b8 = 16'b1110111100100110;
wire v4b9 = v4b8 == v9b;
wire v4ba = v4b9 & ved & v2d0;
wire v4bb = v8b & v22 & v25 & v8f & v31 & v34 & v37 & v3a & vdb & v42 & v45 & v48 & v4a & v4d & v50 & v53 & v477 & v5b & v478 & v60 & v63 & v66;
wire v4bc = v4b7 & v13 & v8a & v11 & v2d2 & v2d3 & v119 & v4ba & v78 & v4bb & v7a & vf0 & v2d4 & v2d5 & v4b0 & v4b1;
wire rnx2x95 = rnx2x94 || v4bc;
wire onx2x95 = onx2x94 || ( rnx2x94 && v4bc);
wire [15:0] v4bd = 16'b1110111100100100;
wire v4be = v4bd == v9b;
wire v4bf = v143;
wire v4c0 = v4bf ^ v72;
wire v4c1 = v4c0 & v72 & v493;
wire v4c2 = v4be & v21f & v115 & v4c1;
wire v4c3 = v484 & v11 & v42f & v13 & v8a & v2d2 & v119 & v78 & v4c2 & v7a & vf0 & v2d5 & v4b0 & v4b1;
wire rnx2x96 = rnx2x95 || v4c3;
wire onx2x96 = onx2x95 || ( rnx2x95 && v4c3);
wire v4c4 = v4b9 & v4a1 & ved & v73;
wire v4c5 = v4bb & v44d & v11 & v2d2 & v119 & v13 & v4c4 & v8a & v78 & v7a & vf0 & v2d5 & v4b0 & v4b1;
wire rnx2x97 = rnx2x96 || v4c5;
wire onx2x97 = onx2x96 || ( rnx2x96 && v4c5);
wire v4c6 = v8b & v22 & v25 & v8f & v31 & v34 & v37 & v3a & v3f & v42 & v45 & v48 & v4a & v4d & v50 & v53 & v477 & v5b & v478 & v60 & v63 & v66;
wire v4c7 = v266 == Advice_1;
wire [23:0] v4c8 = 24'b011001001110111100100101;
wire v4c9 = v4c8 == vaf;
wire v4ca = v4c9 & v71 & v2d0;
wire v4cb = v4c6 & v4c7 & v11 & v8a & v453 & v13 & v428 & v4ca & v78 & ve0 & v7a & vf0 & v2d4 & v401 & v4b0 & v4b1;
wire rnx2x98 = rnx2x97 || v4cb;
wire onx2x98 = onx2x97 || ( rnx2x97 && v4cb);
wire v4cc = v8b & v22 & v25 & v8f & v31 & v34 & v37 & v3a & v170 & v42 & v45 & v48 & v4a & v4d & v50 & v53 & v477 & v5b & v478 & v60 & v63 & v66;
wire [23:0] v4cd = 24'b101001101110111100100110;
wire v4ce = v4cd == vaf;
wire v4cf = v4ce & v16c & v2d0;
wire [31:0] v4d0 = v3e5 + v174;
wire v4d1 = v4d0 == Advice_1;
wire v4d2 = Advice_13 == Advice_30;
wire v4d3 = v4cc & v8a & v11 & v453 & v428 & v13 & ve0 & v4cf & v78 & v4d1 & v7a & vf0 & v2d4 & v4d2 & v4b0 & v4b1;
wire rnx2x99 = rnx2x98 || v4d3;
wire onx2x99 = onx2x98 || ( rnx2x98 && v4d3);
wire v2 = (!onx2x99) && rnx2x99;
assign result = v2;
assign dummy = 1'b0;
endmodule
