module circuit(
input [1544:0] current,
input [1544:0] next,

output [0:0] result,
output [0:0] dummy
);
wire [31:0] Advice_1 = current[31: 0];
wire [1:0] Advice_10 = current[33: 32];
wire [1:0] Advice_11 = current[35: 34];
wire [1:0] Advice_12 = current[37: 36];
wire [1:0] Advice_13 = current[39: 38];
wire [1:0] Advice_14 = current[41: 40];
wire Advice_15 = current[42: 42];
wire Advice_16 = current[43: 43];
wire Advice_17 = current[44: 44];
wire [2:0] Advice_18 = current[47: 45];
wire Advice_19 = current[48: 48];
wire [2:0] Advice_2 = current[51: 49];
wire [2:0] Advice_20 = current[54: 52];
wire Advice_21 = current[55: 55];
wire [2:0] Advice_22 = current[58: 56];
wire Advice_23 = current[59: 59];
wire [31:0] Advice_24 = current[91: 60];
wire [2:0] Advice_25 = current[94: 92];
wire [31:0] Advice_26 = current[126: 95];
wire [2:0] Advice_27 = current[129: 127];
wire Advice_28 = current[130: 130];
wire [2:0] Advice_29 = current[133: 131];
wire [2:0] Advice_3 = current[136: 134];
wire [2:0] Advice_30 = current[139: 137];
wire [1:0] Advice_31 = current[141: 140];
wire [2:0] Advice_32 = current[144: 142];
wire [2:0] Advice_4 = current[147: 145];
wire [2:0] Advice_5 = current[150: 148];
wire [2:0] Advice_6 = current[153: 151];
wire [2:0] Advice_7 = current[156: 154];
wire [2:0] Advice_8 = current[159: 157];
wire [2:0] Advice_9 = current[162: 160];
wire In_error_flag = current[163: 163];
wire In_register_AF = current[428: 428];
wire In_register_CF = current[429: 429];
wire [31:0] In_register_CSBASE = current[461: 430];
wire [7:0] In_register_DF = current[469: 462];
wire [31:0] In_register_DSBASE = current[501: 470];
wire [31:0] In_register_EAX = current[533: 502];
wire [31:0] In_register_EBP = current[565: 534];
wire [31:0] In_register_EBX = current[597: 566];
wire [31:0] In_register_ECX = current[629: 598];
wire [31:0] In_register_EDI = current[661: 630];
wire [31:0] In_register_EDX = current[693: 662];
wire [31:0] In_register_EIP = current[725: 694];
wire [31:0] In_register_ESBASE = current[757: 726];
wire [31:0] In_register_ESI = current[789: 758];
wire [31:0] In_register_ESP = current[821: 790];
wire [31:0] In_register_FSBASE = current[853: 822];
wire [31:0] In_register_GSBASE = current[885: 854];
wire In_register_OF = current[886: 886];
wire In_register_PF = current[887: 887];
wire In_register_SF = current[888: 888];
wire [31:0] In_register_SSBASE = current[920: 889];
wire In_register_ZF = current[921: 921];
wire [63:0] In_timestamp = current[985: 922];
wire Out_error_flag = next[163: 163];
wire Out_register_AF = next[428: 428];
wire Out_register_CF = next[429: 429];
wire [31:0] Out_register_CSBASE = next[461: 430];
wire [7:0] Out_register_DF = next[469: 462];
wire [31:0] Out_register_DSBASE = next[501: 470];
wire [31:0] Out_register_EAX = next[533: 502];
wire [31:0] Out_register_EBP = next[565: 534];
wire [31:0] Out_register_EBX = next[597: 566];
wire [31:0] Out_register_ECX = next[629: 598];
wire [31:0] Out_register_EDI = next[661: 630];
wire [31:0] Out_register_EDX = next[693: 662];
wire [31:0] Out_register_EIP = next[725: 694];
wire [31:0] Out_register_ESBASE = next[757: 726];
wire [31:0] Out_register_ESI = next[789: 758];
wire [31:0] Out_register_ESP = next[821: 790];
wire [31:0] Out_register_FSBASE = next[853: 822];
wire [31:0] Out_register_GSBASE = next[885: 854];
wire Out_register_OF = next[886: 886];
wire Out_register_PF = next[887: 887];
wire Out_register_SF = next[888: 888];
wire [31:0] Out_register_SSBASE = next[920: 889];
wire Out_register_ZF = next[921: 921];
wire [63:0] Out_timestamp = next[985: 922];
wire [119:0] instruction_bits = current[283: 164];
wire [143:0] memory_0 = current[427: 284];
wire v2f = 1'b0;
wire v31 = v2f == Out_error_flag;
wire v33 = In_error_flag == v2f;
wire [3:0] v35 = 4'b0010;
wire v38 =  v35 == memory_0[15: 12] && Advice_1 == memory_0[47: 16] && In_timestamp == memory_0[143: 80] && 4'd0 == memory_0[11: 8] && 1'b1 == memory_0[0: 0] && 6'b000000 == memory_0[7: 2] && 1'b0 == memory_0[1: 1];
wire [2:0] v39 = instruction_bits[29: 27];
wire [2:0] v3a = { v39 };
wire v3c = v3a == Advice_2;
wire [31:0] v3d = memory_0[79: 48];
wire [63:0] v3e = { 32'b00000000000000000000000000000000, v3d };
wire [63:0] v3f = { 32'b00000000000000000000000000000000, In_register_EAX };
wire [63:0] v40 = v3e * v3f;
wire [31:0] v41 = v40[31:0];
wire v42 = v41 == Out_register_EAX;
wire v43 = In_register_EBX == Out_register_EBX;
wire v44 = In_register_ECX == Out_register_ECX;
wire [63:0] v45 = 64'b0000010000000000000000000000000000000000000000000000000000000000;
wire [63:0] v46 = v40 >> v45;
wire [31:0] v47 = v46[31:0];
wire v48 = v47 == Out_register_EDX;
wire v49 = In_register_ESI == Out_register_ESI;
wire v4a = In_register_EDI == Out_register_EDI;
wire v4b = In_register_ESP == Out_register_ESP;
wire v4c = In_register_EBP == Out_register_EBP;
wire [31:0] v4d = 32'b10100000000000000000000000000000;
wire [31:0] v4e = In_register_EIP + v4d;
wire v4f = v4e == Out_register_EIP;
wire v50 = In_register_CSBASE == Out_register_CSBASE;
wire v51 = In_register_SSBASE == Out_register_SSBASE;
wire v52 = In_register_ESBASE == Out_register_ESBASE;
wire v53 = In_register_DSBASE == Out_register_DSBASE;
wire v54 = In_register_GSBASE == Out_register_GSBASE;
wire v55 = In_register_FSBASE == Out_register_FSBASE;
wire v56 = In_register_AF == Out_register_AF;
wire [63:0] v57 = 64'b1111111111111111111111111111111100000000000000000000000000000000;
wire v58 = v40 > v57;
wire v59 = v58 == Out_register_CF;
wire v5a = In_register_DF == Out_register_DF;
wire v5b = v58 == Out_register_OF;
wire v5c = In_register_PF == Out_register_PF;
wire v5d = In_register_SF == Out_register_SF;
wire v5e = In_register_ZF == Out_register_ZF;
wire v5f = v42 & v43 & v44 & v48 & v49 & v4a & v4b & v4c & v4f & v50 & v51 & v52 & v53 & v54 & v55 & v56 & v59 & v5a & v5b & v5c & v5d & v5e;
wire [23:0] v60 = 24'b101001101110111100100110;
wire [23:0] v61 = instruction_bits[23: 0];
wire v62 = v60 == v61;
wire [79:0] v63 = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
wire [79:0] v64 = instruction_bits[119: 40];
wire v65 = v63 == v64;
wire v66 = 1'b1;
wire [2:0] v67 = 3'b001;
wire v68 = Advice_2 == v67;
wire v69 = v68;
wire v6a = v69 ^ v66;
wire v6b = v66 & v6a & v66;
wire v6c = v62 & v65 & v6b;
wire [63:0] v6d = 64'b1000000000000000000000000000000000000000000000000000000000000000;
wire [63:0] v6e = In_timestamp + v6d;
wire v70 = v6e == Out_timestamp;
wire [31:0] v72 = ( Advice_3 == 3'd0) ? In_register_GSBASE :
	( Advice_3 == 3'd1) ? In_register_GSBASE :
	( Advice_3 == 3'd2) ? In_register_GSBASE :
	( Advice_3 == 3'd3) ? In_register_GSBASE :
	( Advice_3 == 3'd4) ? In_register_GSBASE :
	( Advice_3 == 3'd5) ? In_register_GSBASE :
	( Advice_3 == 3'd6) ? In_register_GSBASE : In_register_GSBASE;
wire [31:0] v74 = ( Advice_4 == 3'd0) ? In_register_EAX :
	( Advice_4 == 3'd1) ? In_register_ECX :
	( Advice_4 == 3'd2) ? In_register_EDX :
	( Advice_4 == 3'd3) ? In_register_EBX :
	( Advice_4 == 3'd4) ? In_register_ESP :
	( Advice_4 == 3'd5) ? In_register_EBP :
	( Advice_4 == 3'd6) ? In_register_ESI : In_register_EDI;
wire [31:0] v75 = v72 + v74;
wire [31:0] v77 = ( Advice_5 == 3'd0) ? In_register_EAX :
	( Advice_5 == 3'd1) ? In_register_ECX :
	( Advice_5 == 3'd2) ? In_register_EDX :
	( Advice_5 == 3'd3) ? In_register_EBX :
	( Advice_5 == 3'd4) ? In_register_ESP :
	( Advice_5 == 3'd5) ? In_register_EBP :
	( Advice_5 == 3'd6) ? In_register_ESI : In_register_EDI;
wire [1:0] v78 = instruction_bits[31: 30];
wire [31:0] v79 = { 30'b000000000000000000000000000000, v78 };
wire [31:0] v7b = v77 << v79;
wire [31:0] v7c = v75 + v7b;
wire [7:0] v7d = instruction_bits[39: 32];
wire [7:0] pad_126 = (v7d[7:7] == 1'b1) ?24'b111111111111111111111111 : 24'b000000000000000000000000;
wire [31:0] v7e = { pad_126, v7d };
wire [31:0] v80 = v7c + v7e;
wire v81 = v80 == Advice_1;
wire [2:0] v82 = instruction_bits[26: 24];
wire [2:0] v83 = { v82 };
wire v85 = v83 == Advice_6;
wire v87 = v83 == Advice_7;
wire v88 = In_error_flag ^ v66;
wire v89 = v88 | Out_error_flag;
wire v8a = Advice_6 == Advice_4;
wire v8b = Advice_2 == Advice_5;
wire v8c = Advice_7 == Advice_3;
wire v8d = v31 & v33 & v38 & v3c & v5f & v6c & v70 & v81 & v85 & v87 & v89 & v8a & v8b & v8c;
wire rnx46x0 = 1'b0 || v8d;
wire onx46x0 = 1'b0 || ( 1'b0 && v8d);
wire [31:0] v8e = 32'b00010000000000000000000000000000;
wire [31:0] v8f = In_register_EIP + v8e;
wire v90 = v8f == Out_register_EIP;
wire v91 = v42 & v43 & v44 & v48 & v49 & v4a & v4b & v4c & v90 & v50 & v51 & v52 & v53 & v54 & v55 & v56 & v59 & v5a & v5b & v5c & v5d & v5e;
wire [31:0] v93 = ( Advice_8 == 3'd0) ? In_register_ESBASE :
	( Advice_8 == 3'd1) ? In_register_ESBASE :
	( Advice_8 == 3'd2) ? In_register_ESBASE :
	( Advice_8 == 3'd3) ? In_register_ESBASE :
	( Advice_8 == 3'd4) ? In_register_ESBASE :
	( Advice_8 == 3'd5) ? In_register_ESBASE :
	( Advice_8 == 3'd6) ? In_register_ESBASE : In_register_ESBASE;
wire [31:0] v94 = v93 + v74;
wire [31:0] v95 = v94 + v7b;
wire [31:0] v96 = instruction_bits[63: 32];
wire [31:0] v98 = v95 + v96;
wire v99 = v98 == Advice_1;
wire [23:0] v9a = 24'b011001001110111100100101;
wire v9b = v9a == v61;
wire [55:0] v9c = 56'b00000000000000000000000000000000000000000000000000000000;
wire [55:0] v9d = instruction_bits[119: 64];
wire v9e = v9c == v9d;
wire v9f = v9b & v9e & v6b;
wire va0 = Advice_7 == Advice_8;
wire va1 = v31 & v33 & v91 & v99 & v3c & v85 & v70 & v9f & v38 & v87 & v89 & v8a & v8b & va0;
wire rnx46x1 = rnx46x0 || va1;
wire onx46x1 = onx46x0 || ( rnx46x0 && va1);
wire [31:0] va2 = 32'b00100000000000000000000000000000;
wire [31:0] va3 = In_register_EIP + va2;
wire va4 = va3 == Out_register_EIP;
wire va5 = v42 & v43 & v44 & v48 & v49 & v4a & v4b & v4c & va4 & v50 & v51 & v52 & v53 & v54 & v55 & v56 & v59 & v5a & v5b & v5c & v5d & v5e;
wire [31:0] va7 = ( Advice_9 == 3'd0) ? In_register_DSBASE :
	( Advice_9 == 3'd1) ? In_register_DSBASE :
	( Advice_9 == 3'd2) ? In_register_DSBASE :
	( Advice_9 == 3'd3) ? In_register_DSBASE :
	( Advice_9 == 3'd4) ? In_register_SSBASE :
	( Advice_9 == 3'd5) ? In_register_SSBASE :
	( Advice_9 == 3'd6) ? In_register_DSBASE : In_register_DSBASE;
wire [31:0] va8 = va7 + v74;
wire [31:0] va9 = 32'b00000000000000000000000000000000;
wire [31:0] vab = va9 << va9;
wire [31:0] vac = va8 + vab;
wire [7:0] vad = instruction_bits[31: 24];
wire [7:0] pad_174 = (vad[7:7] == 1'b1) ?24'b111111111111111111111111 : 24'b000000000000000000000000;
wire [31:0] vae = { pad_174, vad };
wire [31:0] vb0 = vac + vae;
wire vb1 = vb0 == Advice_1;
wire [2:0] vb2 = instruction_bits[18: 16];
wire [2:0] vb3 = { vb2 };
wire vb4 = vb3 == Advice_7;
wire vb5 = vb3 == Advice_6;
wire [15:0] vb6 = 16'b1110111100100110;
wire [15:0] vb7 = instruction_bits[15: 0];
wire vb8 = vb6 == vb7;
wire [4:0] vb9 = 5'b00101;
wire [4:0] vba = instruction_bits[23: 19];
wire vbb = vb9 == vba;
wire [87:0] vbc = 88'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
wire [87:0] vbd = instruction_bits[119: 32];
wire vbe = vbc == vbd;
wire vbf = Advice_6 == v67;
wire [2:0] vc0 = 3'b101;
wire vc1 = Advice_6 == vc0;
wire vc2 = vbf & vc1;
wire vc3 = vc2 ^ v66;
wire vc4 = vc3 & v66 & v66;
wire vc5 = vb8 & vbb & vbe & vc4;
wire vc6 = Advice_7 == Advice_9;
wire vc7 = va5 & vb1 & v31 & v33 & v38 & vb4 & vb5 & vc5 & v70 & v89 & v8a & vc6;
wire rnx46x2 = rnx46x1 || vc7;
wire onx46x2 = onx46x1 || ( rnx46x1 && vc7);
wire [31:0] vc8 = 32'b11000000000000000000000000000000;
wire [31:0] vc9 = In_register_EIP + vc8;
wire vca = vc9 == Out_register_EIP;
wire vcb = v42 & v43 & v44 & v48 & v49 & v4a & v4b & v4c & vca & v50 & v51 & v52 & v53 & v54 & v55 & v56 & v59 & v5a & v5b & v5c & v5d & v5e;
wire [31:0] vcc = vac + va9;
wire vcd = vcc == Advice_1;
wire [15:0] vce = 16'b1110111100100100;
wire vcf = vce == vb7;
wire [4:0] vd0 = 5'b00111;
wire vd1 = vd0 == vba;
wire [95:0] vd2 = 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
wire [95:0] vd3 = instruction_bits[119: 24];
wire vd4 = vd2 == vd3;
wire vd5 = vc1;
wire vd6 = vd5 ^ v66;
wire vd7 = Advice_7 == vc0;
wire vd8 = vd7;
wire vd9 = vd8 ^ v66;
wire vda = vd6 & v66 & vd9;
wire vdb = vcf & vd1 & vd4 & vda;
wire vdc = vcb & vcd & v33 & v38 & vb4 & vb5 & v31 & vdb & v70 & v89 & v8a & vc6;
wire rnx46x3 = rnx46x2 || vdc;
wire onx46x3 = onx46x2 || ( rnx46x2 && vdc);
wire [1:0] vdd = instruction_bits[23: 22];
wire [31:0] vde = { 30'b000000000000000000000000000000, vdd };
wire [31:0] ve0 = v77 << vde;
wire [31:0] ve1 = va8 + ve0;
wire [31:0] ve2 = ve1 + vae;
wire ve3 = ve2 == Advice_1;
wire [2:0] ve4 = instruction_bits[21: 19];
wire [2:0] ve5 = { ve4 };
wire ve6 = ve5 == Advice_2;
wire ve7 = vc3 & v6a & v66;
wire ve8 = vb8 & vbe & ve7;
wire ve9 = ve3 & v31 & va5 & v38 & vb4 & v89 & ve6 & v33 & vb5 & ve8 & v70 & v8a & v8b & vc6;
wire rnx46x4 = rnx46x3 || ve9;
wire onx46x4 = onx46x3 || ( rnx46x3 && ve9);
wire [31:0] vea = 32'b01000000000000000000000000000000;
wire [31:0] veb = In_register_EIP + vea;
wire vec = veb == Out_register_EIP;
wire ved = v42 & v43 & v44 & v48 & v49 & v4a & v4b & v4c & vec & v50 & v51 & v52 & v53 & v54 & v55 & v56 & v59 & v5a & v5b & v5c & v5d & v5e;
wire [2:0] vee = instruction_bits[10: 8];
wire [2:0] vef = { vee };
wire vf0 = vef == Advice_6;
wire vf1 = vef == Advice_7;
wire [7:0] vf2 = 8'b11101111;
wire [7:0] vf3 = instruction_bits[7: 0];
wire vf4 = vf2 == vf3;
wire [4:0] vf5 = 5'b00100;
wire [4:0] vf6 = instruction_bits[15: 11];
wire vf7 = vf5 == vf6;
wire [103:0] vf8 = 104'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
wire [103:0] vf9 = instruction_bits[119: 16];
wire vfa = vf8 == vf9;
wire vfb = Advice_7 == v67;
wire vfc = vfb & vd7;
wire vfd = vfc ^ v66;
wire vfe = vc3 & v66 & vfd;
wire vff = vf4 & vf7 & vfa & vfe;
wire v100 = ved & vcd & v31 & v33 & v38 & vf0 & v70 & vf1 & vff & v89 & v8a & vc6;
wire rnx46x5 = rnx46x4 || v100;
wire onx46x5 = onx46x4 || ( rnx46x4 && v100);
wire v101 = instruction_bits[9: 9];
wire v102 = v66 == v101;
wire [4:0] v103 = 5'b00110;
wire v104 = v103 == vf6;
wire v105 = v66 & v66 & v66;
wire v106 = vf4 & v102 & v104 & vd4 & v105;
wire v108 = instruction_bits[8: 8];
wire v107 = instruction_bits[10: 10];
wire [1:0] v109 = { v108 , v107 };
wire v10b = v109 == Advice_10;
wire [31:0] v10d = ( Advice_11 == 2'd0) ? In_register_DSBASE :
	( Advice_11 == 2'd1) ? In_register_DSBASE :
	( Advice_11 == 2'd2) ? In_register_DSBASE : In_register_DSBASE;
wire [31:0] v10f = ( Advice_12 == 2'd0) ? In_register_EDX :
	( Advice_12 == 2'd1) ? In_register_ESI :
	( Advice_12 == 2'd2) ? In_register_EBX : In_register_EDI;
wire [31:0] v110 = v10d + v10f;
wire [31:0] v111 = v110 + vab;
wire [7:0] v112 = instruction_bits[23: 16];
wire [7:0] pad_275 = (v112[7:7] == 1'b1) ?24'b111111111111111111111111 : 24'b000000000000000000000000;
wire [31:0] v113 = { pad_275, v112 };
wire [31:0] v115 = v111 + v113;
wire v116 = v115 == Advice_1;
wire v118 = v109 == Advice_13;
wire v119 = Advice_10 == Advice_12;
wire v11a = Advice_13 == Advice_11;
wire v11b = v33 & v106 & v10b & v116 & v70 & v38 & v118 & vcb & v31 & v89 & v119 & v11a;
wire rnx46x6 = rnx46x5 || v11b;
wire onx46x6 = onx46x5 || ( rnx46x5 && v11b);
wire [31:0] v11c = v74 << v79;
wire [31:0] v11d = v110 + v11c;
wire [31:0] v11e = v11d + va9;
wire v11f = v11e == Advice_1;
wire [31:0] v120 = 32'b00000000111111111111111111111111;
wire [31:0] v121 = In_register_EAX & v120;
wire [7:0] v122 = v3d[7:0];
wire [15:0] v123 = { 8'b00000000, v122 };
wire [7:0] v124 = In_register_EAX[7:0];
wire [15:0] v125 = { 8'b00000000, v124 };
wire [15:0] v126 = v123 * v125;
wire [7:0] v127 = v126[7:0];
wire [31:0] v128 = { 24'b000000000000000000000000, v127 };
wire [31:0] v129 = v121 | v128;
wire [31:0] v12a = 32'b11111111000000001111111111111111;
wire [31:0] v12b = v129 & v12a;
wire [15:0] v12c = 16'b0001000000000000;
wire [15:0] v12d = v126 >> v12c;
wire [7:0] v12e = v12d[7:0];
wire [31:0] v12f = { 24'b000000000000000000000000, v12e };
wire [31:0] v130 = v12f << v8e;
wire [31:0] v131 = v12b | v130;
wire v132 = v131 == Out_register_EAX;
wire v133 = In_register_EDX == Out_register_EDX;
wire [15:0] v134 = 16'b1111111100000000;
wire v135 = v126 > v134;
wire v136 = v135 == Out_register_CF;
wire v137 = v135 == Out_register_OF;
wire v138 = v132 & v43 & v44 & v133 & v49 & v4a & v4b & v4c & va4 & v50 & v51 & v52 & v53 & v54 & v55 & v56 & v136 & v5a & v137 & v5c & v5d & v5e;
wire v13a = instruction_bits[24: 24];
wire v139 = instruction_bits[26: 26];
wire [1:0] v13b = { v13a , v139 };
wire v13c = v13b == Advice_13;
wire v13d = v13b == Advice_10;
wire [23:0] v13e = 24'b011001100110111100100100;
wire v13f = v13e == v61;
wire v140 = instruction_bits[25: 25];
wire v141 = v66 == v140;
wire v142 = v13f & v141 & vbe & v6b;
wire [3:0] v143 = 4'b1000;
wire v144 =  v143 == memory_0[15: 12] && Advice_1 == memory_0[47: 16] && In_timestamp == memory_0[143: 80] && 4'd0 == memory_0[11: 8] && 1'b1 == memory_0[0: 0] && 6'b000000 == memory_0[7: 2] && 1'b0 == memory_0[1: 1];
wire v145 = Advice_2 == Advice_4;
wire v146 = v11f & v138 & v33 & v13c & v13d & v142 & v3c & v70 & v31 & v144 & v89 & v119 & v145 & v11a;
wire rnx46x7 = rnx46x6 || v146;
wire onx46x7 = onx46x6 || ( rnx46x6 && v146);
wire [31:0] v147 = In_register_DSBASE + va9;
wire [31:0] v148 = v74 << vde;
wire [31:0] v149 = v147 + v148;
wire [31:0] v14a = instruction_bits[55: 24];
wire [31:0] v14c = v149 + v14a;
wire v14d = v14c == Advice_1;
wire [31:0] v14e = 32'b11100000000000000000000000000000;
wire [31:0] v14f = In_register_EIP + v14e;
wire v150 = v14f == Out_register_EIP;
wire v151 = v132 & v43 & v44 & v133 & v49 & v4a & v4b & v4c & v150 & v50 & v51 & v52 & v53 & v54 & v55 & v56 & v136 & v5a & v137 & v5c & v5d & v5e;
wire [18:0] v152 = 19'b0110111100100100101;
wire [18:0] v153 = instruction_bits[18: 0];
wire v154 = v152 == v153;
wire [63:0] v155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
wire [63:0] v156 = instruction_bits[119: 56];
wire v157 = v155 == v156;
wire v158 = v154 & v157 & v6b;
wire v159 = v33 & v14d & v144 & ve6 & v151 & v31 & v158 & v70 & v89 & v145;
wire rnx46x8 = rnx46x7 || v159;
wire onx46x8 = onx46x7 || ( rnx46x7 && v159);
wire [31:0] v15a = vac + v14a;
wire v15b = v15a == Advice_1;
wire [15:0] v15c = 16'b0110011001101111;
wire v15d = v15c == vb7;
wire v15e = vbf;
wire v15f = v15e ^ v66;
wire v160 = vfb;
wire v161 = v160 ^ v66;
wire v162 = v15f & v66 & v161;
wire v163 = v15d & vbb & v157 & v162;
wire v164 = v151 & v15b & v33 & v31 & v144 & vb5 & v163 & vb4 & v70 & v89 & v8a & vc6;
wire rnx46x9 = rnx46x8 || v164;
wire onx46x9 = onx46x8 || ( rnx46x8 && v164);
wire [15:0] v165 = 16'b0110111100100101;
wire v166 = v165 == vb7;
wire v167 = instruction_bits[20: 20];
wire v168 = v66 == v167;
wire v169 = v166 & v168 & v157 & vc4;
wire v16b = instruction_bits[19: 19];
wire v16a = instruction_bits[21: 21];
wire [1:0] v16c = { v16b , v16a };
wire v16e = v16c == Advice_14;
wire [31:0] v16f = v10f << vde;
wire [31:0] v170 = va8 + v16f;
wire [31:0] v171 = v170 + v14a;
wire v172 = v171 == Advice_1;
wire v173 = Advice_14 == Advice_12;
wire v174 = v151 & v31 & v33 & vb4 & v169 & v144 & v16e & v70 & v172 & vb5 & v89 & v8a & v173 & vc6;
wire rnx46x10 = rnx46x9 || v174;
wire onx46x10 = onx46x9 || ( rnx46x9 && v174);
wire v175 = v132 & v43 & v44 & v133 & v49 & v4a & v4b & v4c & vca & v50 & v51 & v52 & v53 & v54 & v55 & v56 & v136 & v5a & v137 & v5c & v5d & v5e;
wire [31:0] v176 = v170 + va9;
wire v177 = v176 == Advice_1;
wire [15:0] v178 = 16'b0110111100100100;
wire v179 = v178 == vb7;
wire v17a = vc3 & v66 & vd9;
wire v17b = v179 & v168 & vd4 & v17a;
wire v17c = v175 & v177 & v144 & v33 & vb4 & v31 & v17b & v16e & vb5 & v70 & v89 & v8a & v173 & vc6;
wire rnx46x11 = rnx46x10 || v17c;
wire onx46x11 = onx46x10 || ( rnx46x10 && v17c);
wire [31:0] v17d = instruction_bits[47: 16];
wire [31:0] v17f = vac + v17d;
wire v180 = v17f == Advice_1;
wire [31:0] v181 = 32'b01100000000000000000000000000000;
wire [31:0] v182 = In_register_EIP + v181;
wire v183 = v182 == Out_register_EIP;
wire v184 = v132 & v43 & v44 & v133 & v49 & v4a & v4b & v4c & v183 & v50 & v51 & v52 & v53 & v54 & v55 & v56 & v136 & v5a & v137 & v5c & v5d & v5e;
wire [7:0] v185 = 8'b01101111;
wire v186 = v185 == vf3;
wire v187 = vb9 == vf6;
wire [71:0] v188 = 72'b000000000000000000000000000000000000000000000000000000000000000000000000;
wire [71:0] v189 = instruction_bits[119: 48];
wire v18a = v188 == v189;
wire v18b = vc3 & v66 & v161;
wire v18c = v186 & v187 & v18a & v18b;
wire v18d = v180 & v184 & v33 & v31 & vf1 & v70 & v144 & vf0 & v18c & v89 & v8a & vc6;
wire rnx46x12 = rnx46x11 || v18d;
wire onx46x12 = onx46x11 || ( rnx46x11 && v18d);
wire [63:0] v18e = { 32'b00000000000000000000000000000000, Advice_1 };
wire [63:0] v18f = v3f * v18e;
wire [31:0] v190 = v18f[31:0];
wire v191 = v190 == Out_register_EAX;
wire [63:0] v192 = v18f >> v45;
wire [31:0] v193 = v192[31:0];
wire v194 = v193 == Out_register_EDX;
wire v195 = v18f > v57;
wire v196 = v195 == Out_register_CF;
wire v197 = v195 == Out_register_OF;
wire v198 = v191 & v43 & v44 & v194 & v49 & v4a & v4b & v4c & vca & v50 & v51 & v52 & v53 & v54 & v55 & v56 & v196 & v5a & v197 & v5c & v5d & v5e;
wire v199 = v74 == Advice_1;
wire [15:0] v19a = 16'b0110110011101111;
wire v19b = v19a == vb7;
wire v19c = v66;
wire v19d = v19b & vd1 & vd4 & v19c;
wire v19e = v198 & v33 & v199 & v89 & v19d & v31 & v70 & vb5 & v8a;
wire rnx46x13 = rnx46x12 || v19e;
wire onx46x13 = onx46x12 || ( rnx46x12 && v19e);
wire v19f = v191 & v43 & v44 & v194 & v49 & v4a & v4b & v4c & vec & v50 & v51 & v52 & v53 & v54 & v55 & v56 & v196 & v5a & v197 & v5c & v5d & v5e;
wire v1a0 = vd0 == vf6;
wire v1a1 = vf4 & v1a0 & vfa & v19c;
wire v1a2 = v19f & v199 & v70 & v33 & vf0 & v31 & v1a1 & v89 & v8a;
wire rnx46x14 = rnx46x13 || v1a2;
wire onx46x14 = onx46x13 || ( rnx46x13 && v1a2);
wire [31:0] v1a4 = ( Advice_15 == 1'd0) ? In_register_EDI : In_register_EBX;
wire [31:0] v1a5 = 32'b11111111111111110000000000000000;
wire [31:0] v1a6 = v1a4 & v1a5;
wire [31:0] v1a7 = v10d + v1a6;
wire [31:0] v1a8 = v1a7 + vab;
wire [31:0] v1a9 = v1a8 + va9;
wire [15:0] v1aa = v1a9[15:0];
wire [31:0] v1ab = { 16'b0000000000000000, v1aa };
wire v1ac = v1ab == Advice_1;
wire [31:0] pad_429 = (v3d[31:31] == 1'b1) ?32'b11111111111111111111111111111111 : 32'b00000000000000000000000000000000;
wire [63:0] v1ad = { pad_429, v3d };
wire [31:0] pad_430 = (In_register_EAX[31:31] == 1'b1) ?32'b11111111111111111111111111111111 : 32'b00000000000000000000000000000000;
wire [63:0] v1ae = { pad_430, In_register_EAX };
wire [63:0] v1af = v1ad * v1ae;
wire [31:0] v1b0 = v1af[31:0];
wire v1b1 = v1b0 == Out_register_EAX;
wire [63:0] v1b2 = v1af >> v45;
wire [31:0] v1b3 = v1b2[31:0];
wire v1b4 = v1b3 == Out_register_EDX;
wire [63:0] v1b5 = 64'b0000000000000000000000000000000111111111111111111111111111111111;
wire [63:0] v1b6 = v1af + v1b5;
wire [63:0] v1b7 = 64'b0000000000000000000000000000000011111111111111111111111111111111;
wire v1b8 = v1b6 < v1b7;
wire v1b9 = v1b8 == Out_register_CF;
wire v1ba = v1b8 == Out_register_OF;
wire v1bb = v1b1 & v43 & v44 & v1b4 & v49 & v4a & v4b & v4c & vca & v50 & v51 & v52 & v53 & v54 & v55 & v56 & v1b9 & v5a & v1ba & v5c & v5d & v5e;
wire v1bc = instruction_bits[17: 17];
wire v1bd = { v1bc };
wire v1bf = v1bd == Advice_16;
wire [16:0] v1c0 = 17'b11100110111011111;
wire [16:0] v1c1 = instruction_bits[16: 0];
wire v1c2 = v1c0 == v1c1;
wire [5:0] v1c3 = 6'b110100;
wire [5:0] v1c4 = instruction_bits[23: 18];
wire v1c5 = v1c3 == v1c4;
wire v1c6 = v1c2 & v1c5 & vd4 & v105;
wire v1c8 = v1bd == Advice_17;
wire v1c9 = Advice_16 == Advice_15;
wire [1:0] v1ca = { Advice_17 , v2f };
wire v1cb = v1ca == Advice_11;
wire v1cc = v1ac & v1bb & v31 & v33 & v38 & v89 & v1bf & v1c6 & v1c8 & v70 & v1c9 & v1cb;
wire rnx46x15 = rnx46x14 || v1cc;
wire onx46x15 = onx46x14 || ( rnx46x14 && v1cc);
wire v1cd = v1b1 & v43 & v44 & v1b4 & v49 & v4a & v4b & v4c & v4f & v50 & v51 & v52 & v53 & v54 & v55 & v56 & v1b9 & v5a & v1ba & v5c & v5d & v5e;
wire [31:0] v1cf = ( Advice_18 == 3'd0) ? In_register_SSBASE :
	( Advice_18 == 3'd1) ? In_register_SSBASE :
	( Advice_18 == 3'd2) ? In_register_SSBASE :
	( Advice_18 == 3'd3) ? In_register_SSBASE :
	( Advice_18 == 3'd4) ? In_register_SSBASE :
	( Advice_18 == 3'd5) ? In_register_SSBASE :
	( Advice_18 == 3'd6) ? In_register_SSBASE : In_register_SSBASE;
wire [31:0] v1d0 = v1cf + v74;
wire [31:0] v1d1 = v1d0 + v7b;
wire [31:0] v1d2 = v1d1 + v7e;
wire v1d3 = v1d2 == Advice_1;
wire [23:0] v1d4 = 24'b011011001110111100110110;
wire v1d5 = v1d4 == v61;
wire v1d6 = v1d5 & v65 & v6b;
wire v1d7 = Advice_7 == Advice_18;
wire v1d8 = v1cd & v33 & v38 & v1d3 & v87 & v1d6 & v85 & v70 & v31 & v3c & v89 & v8a & v8b & v1d7;
wire rnx46x16 = rnx46x15 || v1d8;
wire onx46x16 = onx46x15 || ( rnx46x15 && v1d8);
wire v1d9 = instruction_bits[16: 16];
wire v1da = { v1d9 };
wire v1dc = v1da == Advice_19;
wire [31:0] v1de = ( Advice_20 == 3'd0) ? In_register_EBX :
	( Advice_20 == 3'd1) ? In_register_EBX :
	( Advice_20 == 3'd2) ? In_register_EBP :
	( Advice_20 == 3'd3) ? In_register_EBP :
	( Advice_20 == 3'd4) ? In_register_ESI :
	( Advice_20 == 3'd5) ? In_register_EDI :
	( Advice_20 == 3'd6) ? In_register_EBP : In_register_EBX;
wire [31:0] v1df = v1de & v1a5;
wire [31:0] v1e0 = va7 + v1df;
wire [31:0] v1e2 = ( Advice_21 == 1'd0) ? In_register_ESI : In_register_EDI;
wire [31:0] v1e3 = v1e2 & v1a5;
wire [31:0] v1e4 = 32'b10000000000000000000000000000000;
wire [31:0] v1e6 = v1e3 << v1e4;
wire [31:0] v1e7 = v1e0 + v1e6;
wire [15:0] v1e8 = instruction_bits[39: 24];
wire [15:0] pad_489 = (v1e8[15:15] == 1'b1) ?16'b1111111111111111 : 16'b0000000000000000;
wire [31:0] v1e9 = { pad_489, v1e8 };
wire [31:0] v1eb = v1e7 + v1e9;
wire [15:0] v1ec = v1eb[15:0];
wire [31:0] v1ed = { 16'b0000000000000000, v1ec };
wire v1ee = v1ed == Advice_1;
wire [15:0] v1ef = 16'b1110011011101111;
wire v1f0 = v1ef == vb7;
wire [5:0] v1f1 = 6'b010101;
wire v1f2 = v1f1 == v1c4;
wire v1f3 = Advice_16;
wire v1f4 = v1f3 ^ v66;
wire v1f5 = v1f4 & v66 & v66;
wire v1f6 = v1f0 & v1f2 & v65 & v1f5;
wire [1:0] v1f7 = 2'b00;
wire [2:0] v1f8 = { Advice_16 , v1f7 };
wire v1f9 = v1f8 == Advice_20;
wire v1fa = Advice_19 == Advice_21;
wire [2:0] v1fb = { Advice_17 , v1f7 };
wire v1fc = v1fb == Advice_9;
wire v1fd = v1cd & v33 & v1c8 & v1dc & v70 & v1ee & v31 & v1bf & v1f6 & v38 & v89 & v1f9 & v1fa & v1fc;
wire rnx46x17 = rnx46x16 || v1fd;
wire onx46x17 = onx46x16 || ( rnx46x16 && v1fd);
wire v1fe = v1b1 & v43 & v44 & v1b4 & v49 & v4a & v4b & v4c & v90 & v50 & v51 & v52 & v53 & v54 & v55 & v56 & v1b9 & v5a & v1ba & v5c & v5d & v5e;
wire [23:0] v1ff = 24'b001001101110111100110101;
wire v200 = v1ff == v61;
wire v201 = v200 & v9e & v6b;
wire [31:0] v203 = ( Advice_22 == 3'd0) ? In_register_FSBASE :
	( Advice_22 == 3'd1) ? In_register_FSBASE :
	( Advice_22 == 3'd2) ? In_register_FSBASE :
	( Advice_22 == 3'd3) ? In_register_FSBASE :
	( Advice_22 == 3'd4) ? In_register_FSBASE :
	( Advice_22 == 3'd5) ? In_register_FSBASE :
	( Advice_22 == 3'd6) ? In_register_FSBASE : In_register_FSBASE;
wire [31:0] v204 = v203 + v74;
wire [31:0] v205 = v204 + v7b;
wire [31:0] v206 = v205 + v96;
wire v207 = v206 == Advice_1;
wire v208 = Advice_7 == Advice_22;
wire v209 = v31 & v38 & v87 & v1fe & v3c & v85 & v201 & v70 & v207 & v33 & v89 & v8a & v8b & v208;
wire rnx46x18 = rnx46x17 || v209;
wire onx46x18 = onx46x17 || ( rnx46x17 && v209);
wire v20a = v1b1 & v43 & v44 & v1b4 & v49 & v4a & v4b & v4c & va4 & v50 & v51 & v52 & v53 & v54 & v55 & v56 & v1b9 & v5a & v1ba & v5c & v5d & v5e;
wire [15:0] v20b = 16'b1110111100110110;
wire v20c = v20b == vb7;
wire v20d = v20c & vd1 & vbe & vc4;
wire v20e = v20a & v31 & v33 & v38 & vb5 & v70 & v20d & vb1 & vb4 & v89 & v8a & vc6;
wire rnx46x19 = rnx46x18 || v20e;
wire onx46x19 = onx46x18 || ( rnx46x18 && v20e);
wire [31:0] v20f = v111 + va9;
wire v210 = v20f == Advice_1;
wire v211 = instruction_bits[18: 18];
wire [1:0] v212 = { v1d9 , v211 };
wire v213 = v212 == Advice_10;
wire v214 = v212 == Advice_13;
wire [15:0] v215 = 16'b1110111100110100;
wire v216 = v215 == vb7;
wire v217 = instruction_bits[17: 17];
wire v218 = v66 == v217;
wire v219 = v216 & v218 & vd1 & vd4 & v105;
wire v21a = v1bb & v31 & v33 & v38 & v210 & v213 & v89 & v214 & v70 & v219 & v119 & v11a;
wire rnx46x20 = rnx46x19 || v21a;
wire onx46x20 = onx46x19 || ( rnx46x19 && v21a);
wire [31:0] v21b = v170 + vae;
wire v21c = v21b == Advice_1;
wire [2:0] v21d = 3'b000;
wire v21e = Advice_6 == v21d;
wire [2:0] v21f = 3'b100;
wire v220 = Advice_6 == v21f;
wire [2:0] v221 = 3'b010;
wire v222 = Advice_6 == v221;
wire [2:0] v223 = 3'b110;
wire v224 = Advice_6 == v223;
wire [2:0] v225 = 3'b011;
wire v226 = Advice_6 == v225;
wire [2:0] v227 = 3'b111;
wire v228 = Advice_6 == v227;
wire v229 = v21e & v220 & v222 & v224 & v226 & v228;
wire v22a = v229 ^ v66;
wire v22b = v22a & v66 & v66;
wire v22c = v20c & v168 & vbe & v22b;
wire v22d = v21c & v31 & v38 & v22c & v20a & v33 & v70 & v16e & vb5 & vb4 & v89 & v8a & v173 & vc6;
wire rnx46x21 = rnx46x20 || v22d;
wire onx46x21 = onx46x20 || ( rnx46x20 && v22d);
wire [4:0] v22e = 5'b10110;
wire v22f = v22e == vf6;
wire v230 = vf4 & v102 & v22f & vd4 & v105;
wire v231 = v116 & v1bb & v33 & v31 & v38 & v118 & v70 & v10b & v230 & v89 & v119 & v11a;
wire rnx46x22 = rnx46x21 || v231;
wire onx46x22 = onx46x21 || ( rnx46x21 && v231);
wire v232 = v1b1 & v43 & v44 & v1b4 & v49 & v4a & v4b & v4c & vec & v50 & v51 & v52 & v53 & v54 & v55 & v56 & v1b9 & v5a & v1ba & v5c & v5d & v5e;
wire [4:0] v233 = 5'b10100;
wire v234 = v233 == vf6;
wire v235 = vf4 & v234 & vfa & vfe;
wire v236 = v232 & vcd & v38 & vf0 & vf1 & v235 & v70 & v31 & v33 & v89 & v8a & vc6;
wire rnx46x23 = rnx46x22 || v236;
wire onx46x23 = onx46x22 || ( rnx46x22 && v236);
wire v237 = v1b1 & v43 & v44 & v1b4 & v49 & v4a & v4b & v4c & v183 & v50 & v51 & v52 & v53 & v54 & v55 & v56 & v1b9 & v5a & v1ba & v5c & v5d & v5e;
wire [4:0] v238 = 5'b10101;
wire v239 = v238 == vf6;
wire v23a = vf4 & v239 & v18a & v162;
wire v23b = v237 & v31 & v33 & v180 & v38 & vf1 & v23a & v70 & vf0 & v89 & v8a & vc6;
wire rnx46x24 = rnx46x23 || v23b;
wire onx46x24 = onx46x23 || ( rnx46x23 && v23b);
wire [31:0] v23c = 32'b00000000000000001111111111111111;
wire [31:0] v23d = In_register_EAX & v23c;
wire [15:0] v23e = v3d[15:0];
wire [15:0] pad_575 = (v23e[15:15] == 1'b1) ?16'b1111111111111111 : 16'b0000000000000000;
wire [31:0] v23f = { pad_575, v23e };
wire [15:0] v240 = In_register_EAX[15:0];
wire [15:0] pad_577 = (v240[15:15] == 1'b1) ?16'b1111111111111111 : 16'b0000000000000000;
wire [31:0] v241 = { pad_577, v240 };
wire [31:0] v242 = v23f * v241;
wire [15:0] v243 = v242[15:0];
wire [31:0] v244 = { 16'b0000000000000000, v243 };
wire [31:0] v245 = v23d | v244;
wire v246 = v245 == Out_register_EAX;
wire [31:0] v247 = In_register_EDX & v23c;
wire [31:0] v248 = 32'b00001000000000000000000000000000;
wire [31:0] v249 = v242 >> v248;
wire [15:0] v24a = v249[15:0];
wire [31:0] v24b = { 16'b0000000000000000, v24a };
wire [31:0] v24c = v247 | v24b;
wire v24d = v24c == Out_register_EDX;
wire [31:0] v24e = 32'b00000000000000011111111111111111;
wire [31:0] v24f = v242 + v24e;
wire v250 = v24f < v23c;
wire v251 = v250 == Out_register_CF;
wire v252 = v250 == Out_register_OF;
wire v253 = v246 & v43 & v44 & v24d & v49 & v4a & v4b & v4c & va4 & v50 & v51 & v52 & v53 & v54 & v55 & v56 & v251 & v5a & v252 & v5c & v5d & v5e;
wire [3:0] v254 = 4'b0100;
wire v255 =  v254 == memory_0[15: 12] && Advice_1 == memory_0[47: 16] && In_timestamp == memory_0[143: 80] && 4'd0 == memory_0[11: 8] && 1'b1 == memory_0[0: 0] && 6'b000000 == memory_0[7: 2] && 1'b0 == memory_0[1: 1];
wire [23:0] v256 = 24'b011001101110111100110100;
wire v257 = v256 == v61;
wire v258 = v257 & v141 & vbe & v6b;
wire v259 = v253 & v31 & v255 & v13d & v13c & v89 & v3c & v33 & v70 & v11f & v258 & v119 & v145 & v11a;
wire rnx46x25 = rnx46x24 || v259;
wire onx46x25 = onx46x24 || ( rnx46x24 && v259);
wire [31:0] v25b = 32'b00000000000000000000000000000000;
wire [31:0] v25c = ( Advice_23 == 1'd0) ? v25b : In_register_EBP;
wire [31:0] v25d = v25c & v1a5;
wire [31:0] v25e = va7 + v25d;
wire [31:0] v25f = v25e + v1e6;
wire [31:0] v260 = v25f + vae;
wire [15:0] v261 = v260[15:0];
wire [31:0] v262 = { 16'b0000000000000000, v261 };
wire v263 = v262 == Advice_1;
wire [15:0] v264 = 16'b1110011001101111;
wire v265 = v264 == vb7;
wire [5:0] v266 = 6'b010110;
wire v267 = v266 == v1c4;
wire v268 = Advice_23 == v2f;
wire v269 = v268;
wire v26a = v269 ^ v66;
wire v26b = v26a & v66 & v66;
wire v26c = v265 & v267 & vbe & v26b;
wire [7:0] pad_621 = (v122[7:7] == 1'b1) ?8'b11111111 : 8'b00000000;
wire [15:0] v26d = { pad_621, v122 };
wire [7:0] pad_622 = (v124[7:7] == 1'b1) ?8'b11111111 : 8'b00000000;
wire [15:0] v26e = { pad_622, v124 };
wire [15:0] v26f = v26d * v26e;
wire [7:0] v270 = v26f[7:0];
wire [31:0] v271 = { 24'b000000000000000000000000, v270 };
wire [31:0] v272 = v121 | v271;
wire [31:0] v273 = v272 & v12a;
wire [15:0] v274 = v26f >> v12c;
wire [7:0] v275 = v274[7:0];
wire [31:0] v276 = { 24'b000000000000000000000000, v275 };
wire [31:0] v277 = v276 << v8e;
wire [31:0] v278 = v273 | v277;
wire v279 = v278 == Out_register_EAX;
wire [15:0] v27a = 16'b0000000111111111;
wire [15:0] v27b = v26f + v27a;
wire [15:0] v27c = 16'b0000000011111111;
wire v27d = v27b < v27c;
wire v27e = v27d == Out_register_CF;
wire v27f = v27d == Out_register_OF;
wire v280 = v279 & v43 & v44 & v133 & v49 & v4a & v4b & v4c & va4 & v50 & v51 & v52 & v53 & v54 & v55 & v56 & v27e & v5a & v27f & v5c & v5d & v5e;
wire v281 = Advice_16 == Advice_23;
wire v282 = v263 & v144 & v31 & v33 & v1c8 & v89 & v26c & v280 & v70 & v1dc & v1bf & v281 & v1fa & v1fc;
wire rnx46x26 = rnx46x25 || v282;
wire onx46x26 = onx46x25 || ( rnx46x25 && v282);
wire v283 = v279 & v43 & v44 & v133 & v49 & v4a & v4b & v4c & vca & v50 & v51 & v52 & v53 & v54 & v55 & v56 & v27e & v5a & v27f & v5c & v5d & v5e;
wire [31:0] v284 = v25f + va9;
wire [15:0] v285 = v284[15:0];
wire [31:0] v286 = { 16'b0000000000000000, v285 };
wire v287 = v286 == Advice_1;
wire [5:0] v288 = 6'b010100;
wire v289 = v288 == v1c4;
wire v28a = v265 & v289 & vd4 & v26b;
wire v28b = v283 & v287 & v144 & v31 & v1c8 & v28a & v1dc & v70 & v33 & v1bf & v89 & v281 & v1fa & v1fc;
wire rnx46x27 = rnx46x26 || v28b;
wire onx46x27 = onx46x26 || ( rnx46x26 && v28b);
wire v28c = v279 & v43 & v44 & v133 & v49 & v4a & v4b & v4c & v150 & v50 & v51 & v52 & v53 & v54 & v55 & v56 & v27e & v5a & v27f & v5c & v5d & v5e;
wire [18:0] v28d = 19'b0110111100110100101;
wire v28e = v28d == v153;
wire v28f = v28e & v157 & v6b;
wire v290 = v33 & v144 & ve6 & v28c & v14d & v28f & v31 & v70 & v89 & v145;
wire rnx46x28 = rnx46x27 || v290;
wire onx46x28 = onx46x27 || ( rnx46x27 && v290);
wire [31:0] v291 = v94 + vab;
wire [31:0] v292 = v291 + v14a;
wire v293 = v292 == Advice_1;
wire [15:0] v294 = 16'b0110010001101111;
wire v295 = v294 == vb7;
wire v296 = v238 == vba;
wire v297 = v295 & v296 & v157 & v162;
wire v298 = v28c & v31 & v33 & v144 & v293 & v89 & vb4 & v70 & vb5 & v297 & v8a & va0;
wire rnx46x29 = rnx46x28 || v298;
wire onx46x29 = onx46x28 || ( rnx46x28 && v298);
wire [31:0] v299 = v110 + v148;
wire [31:0] v29a = v299 + va9;
wire v29b = v29a == Advice_1;
wire [15:0] v29c = 16'b0110111100110100;
wire v29d = v29c == vb7;
wire v29e = v29d & v218 & vd4 & v6b;
wire v29f = v144 & v283 & v214 & v29b & v31 & ve6 & v29e & v213 & v70 & v33 & v89 & v119 & v145 & v11a;
wire rnx46x30 = rnx46x29 || v29f;
wire onx46x30 = onx46x29 || ( rnx46x29 && v29f);
wire v2a1 = v96 == Advice_24;
wire [31:0] pad_674 = (Advice_24[31:31] == 1'b1) ?32'b11111111111111111111111111111111 : 32'b00000000000000000000000000000000;
wire [63:0] v2a2 = { pad_674, Advice_24 };
wire [63:0] v2a3 = v1ad * v2a2;
wire [31:0] v2a4 = v2a3[31:0];
wire [31:0] v2a5 = { v2a4 };
wire [31:0] v2a7 = ( Advice_25 == 3'd0) ? Out_register_EAX :
	( Advice_25 == 3'd1) ? Out_register_ECX :
	( Advice_25 == 3'd2) ? Out_register_EDX :
	( Advice_25 == 3'd3) ? Out_register_EBX :
	( Advice_25 == 3'd4) ? Out_register_ESP :
	( Advice_25 == 3'd5) ? Out_register_EBP :
	( Advice_25 == 3'd6) ? Out_register_ESI : Out_register_EDI;
wire v2a8 = v2a5 == v2a7;
wire v2a9 = In_register_EAX == Out_register_EAX;
wire v2aa = v21e | v2a9;
wire v2ab = v224 | v43;
wire v2ac = v220 | v44;
wire v2ad = v222 | v133;
wire v2ae = v226 | v49;
wire v2af = v228 | v4a;
wire v2b0 = vbf | v4b;
wire v2b1 = vc1 | v4c;
wire [63:0] v2b2 = v2a3 + v1b5;
wire v2b3 = v2b2 < v1b7;
wire v2b4 = v2b3 == Out_register_CF;
wire v2b5 = v2b3 == Out_register_OF;
wire v2b6 = v2aa & v2ab & v2ac & v2ad & v2ae & v2af & v2b0 & v2b1 & v90 & v50 & v51 & v52 & v53 & v54 & v55 & v56 & v2b4 & v5a & v2b5 & v5c & v5d & v5e;
wire v2b7 = v2a8 & v2b6;
wire v2b9 =  v35 == memory_0[15: 12] && Advice_26 == memory_0[47: 16] && In_timestamp == memory_0[143: 80] && 4'd0 == memory_0[11: 8] && 1'b1 == memory_0[0: 0] && 6'b000000 == memory_0[7: 2] && 1'b0 == memory_0[1: 1];
wire v2ba = v3a == Advice_7;
wire v2bc = v83 == Advice_27;
wire v2bd = v83 == Advice_2;
wire [18:0] v2be = 19'b1010011010010110001;
wire v2bf = v2be == v153;
wire v2c0 = v1f7 == vdd;
wire v2c1 = Advice_2 == vc0;
wire v2c2 = v2c1;
wire v2c3 = v2c2 ^ v66;
wire v2c4 = Advice_27 == vc0;
wire v2c5 = v2c4;
wire v2c6 = v2c5 ^ v66;
wire v2c7 = v66 & v2c3 & v161 & v2c6;
wire v2c8 = v2bf & v2c0 & v9e & v2c7;
wire [31:0] v2c9 = v7c + va9;
wire v2ca = v2c9 == Advice_26;
wire v2cb = ve5 == Advice_6;
wire v2cc = Advice_7 == Advice_5;
wire v2cd = Advice_27 == Advice_3;
wire v2ce = Advice_6 == Advice_25;
wire v2cf = v2a1 & v2b7 & v31 & v2b9 & v2ba & v2bc & v2bd & v2c8 & v2ca & v33 & v2cb & v70 & v89 & v145 & v2cc & v2cd & v2ce;
wire rnx46x31 = rnx46x30 || v2cf;
wire onx46x31 = onx46x30 || ( rnx46x30 && v2cf);
wire v2d0 = v14a == Advice_24;
wire v2d1 = v2aa & v2ab & v2ac & v2ad & v2ae & v2af & v2b0 & v2b1 & v150 & v50 & v51 & v52 & v53 & v54 & v55 & v56 & v2b4 & v5a & v2b5 & v5c & v5d & v5e;
wire v2d2 = v2a8 & v2d1;
wire v2d3 = v286 == Advice_26;
wire v2d4 = v1da == Advice_17;
wire [15:0] v2d5 = 16'b1110011010010110;
wire v2d6 = v2d5 == vb7;
wire v2d7 = instruction_bits[18: 18];
wire v2d8 = v2f == v2d7;
wire v2d9 = v66 & v26a & v66 & v66;
wire v2da = v2d6 & v2d8 & v2c0 & v157 & v2d9;
wire v2db = v1bd == Advice_19;
wire v2dd = v1bd == Advice_28;
wire v2de = Advice_19 == Advice_23;
wire v2df = Advice_17 == Advice_21;
wire [2:0] v2e0 = { Advice_28 , v1f7 };
wire v2e1 = v2e0 == Advice_9;
wire v2e2 = v2d0 & v2d2 & v70 & v2d3 & v31 & v33 & v2b9 & v2d4 & v2da & v2db & v2cb & v2dd & v89 & v2de & v2df & v2e1 & v2ce;
wire rnx46x32 = rnx46x31 || v2e2;
wire onx46x32 = onx46x31 || ( rnx46x31 && v2e2);
wire [31:0] v2e3 = v10d + v1e3;
wire [31:0] v2e4 = v2e3 + vab;
wire [31:0] v2e5 = v2e4 + va9;
wire [15:0] v2e6 = v2e5[15:0];
wire [31:0] v2e7 = { 16'b0000000000000000, v2e6 };
wire v2e8 = v2e7 == Advice_26;
wire v2e9 = v1da == Advice_28;
wire [1:0] v2ea = 2'b01;
wire [1:0] v2eb = instruction_bits[18: 17];
wire v2ec = v2ea == v2eb;
wire v2ed = v66 & v66 & v66 & v66;
wire v2ee = v2d6 & v2ec & v2c0 & v157 & v2ed;
wire [1:0] v2ef = { Advice_28 , v2f };
wire v2f0 = v2ef == Advice_11;
wire v2f1 = v2d2 & v2d0 & v2cb & v2e8 & v31 & v33 & v70 & v2b9 & v2e9 & v89 & v1dc & v2ee & v1fa & v2f0 & v2ce;
wire rnx46x33 = rnx46x32 || v2f1;
wire onx46x33 = onx46x32 || ( rnx46x32 && v2f1);
wire [31:0] v2f2 = 32'b11010000000000000000000000000000;
wire [31:0] v2f3 = In_register_EIP + v2f2;
wire v2f4 = v2f3 == Out_register_EIP;
wire v2f5 = v2aa & v2ab & v2ac & v2ad & v2ae & v2af & v2b0 & v2b1 & v2f4 & v50 & v51 & v52 & v53 & v54 & v55 & v56 & v2b4 & v5a & v2b5 & v5c & v5d & v5e;
wire v2f6 = v2a8 & v2f5;
wire [31:0] v2f7 = instruction_bits[87: 56];
wire v2f9 = v2f7 == Advice_24;
wire [31:0] v2fa = In_register_GSBASE + va9;
wire [31:0] v2fb = v2fa + vab;
wire [31:0] v2fc = v2fb + v14a;
wire v2fd = v2fc == Advice_26;
wire [18:0] v2fe = 19'b1010011010010110101;
wire v2ff = v2fe == v153;
wire [31:0] v300 = instruction_bits[119: 88];
wire v301 = va9 == v300;
wire v302 = v2ff & v2c0 & v301 & v2ed;
wire v303 = v2f6 & v2f9 & v2fd & v31 & v302 & v2b9 & v2cb & v70 & v33 & v89 & v2ce;
wire rnx46x34 = rnx46x33 || v303;
wire onx46x34 = onx46x33 || ( rnx46x33 && v303);
wire [31:0] v304 = 32'b00110000000000000000000000000000;
wire [31:0] v305 = In_register_EIP + v304;
wire v306 = v305 == Out_register_EIP;
wire v307 = v2aa & v2ab & v2ac & v2ad & v2ae & v2af & v2b0 & v2b1 & v306 & v50 & v51 & v52 & v53 & v54 & v55 & v56 & v2b4 & v5a & v2b5 & v5c & v5d & v5e;
wire v308 = v2a8 & v307;
wire [31:0] v309 = instruction_bits[95: 64];
wire v30b = v309 == Advice_24;
wire [31:0] v30c = v1d1 + v96;
wire v30d = v30c == Advice_26;
wire [18:0] v30e = 19'b0110110010010110001;
wire v30f = v30e == v153;
wire v310 = v2ea == vdd;
wire [23:0] v311 = 24'b000000000000000000000000;
wire [23:0] v312 = instruction_bits[119: 96];
wire v313 = v311 == v312;
wire v314 = v66 & v66 & v161 & v66;
wire v315 = v30f & v310 & v313 & v314;
wire v316 = Advice_27 == Advice_18;
wire v317 = v308 & v30b & v2bc & v33 & v31 & v2ba & v2b9 & v2bd & v30d & v2cb & v70 & v315 & v89 & v145 & v2cc & v316 & v2ce;
wire rnx46x35 = rnx46x34 || v317;
wire onx46x35 = onx46x34 || ( rnx46x34 && v317);
wire [31:0] v319 = ( Advice_29 == 3'd0) ? In_register_DSBASE :
	( Advice_29 == 3'd1) ? In_register_DSBASE :
	( Advice_29 == 3'd2) ? In_register_SSBASE :
	( Advice_29 == 3'd3) ? In_register_SSBASE :
	( Advice_29 == 3'd4) ? In_register_DSBASE :
	( Advice_29 == 3'd5) ? In_register_DSBASE :
	( Advice_29 == 3'd6) ? In_register_SSBASE : In_register_DSBASE;
wire [31:0] v31a = v319 + v1df;
wire [31:0] v31c = ( Advice_30 == 3'd0) ? In_register_ESI :
	( Advice_30 == 3'd1) ? In_register_EDI :
	( Advice_30 == 3'd2) ? In_register_ESI :
	( Advice_30 == 3'd3) ? In_register_EDI :
	( Advice_30 == 3'd4) ? va9 :
	( Advice_30 == 3'd5) ? va9 :
	( Advice_30 == 3'd6) ? va9 : va9;
wire [31:0] v31d = v31c & v1a5;
wire [31:0] v31e = v31d << v1e4;
wire [31:0] v31f = v31a + v31e;
wire [31:0] v320 = v31f + vae;
wire [15:0] v321 = v320[15:0];
wire [31:0] v322 = { 16'b0000000000000000, v321 };
wire v323 = v322 == Advice_26;
wire v324 = vb3 == Advice_27;
wire [1:0] v325 = 2'b10;
wire v326 = v325 == vdd;
wire v327 = v2d6 & v326 & v9e & v2ed;
wire v328 = vb3 == Advice_2;
wire v329 = Advice_2 == Advice_20;
wire v32a = Advice_7 == Advice_30;
wire v32b = Advice_27 == Advice_29;
wire v32c = v2a1 & v323 & v31 & v2cb & v2b9 & v324 & v2b7 & vb4 & v327 & v328 & v33 & v70 & v89 & v329 & v32a & v32b & v2ce;
wire rnx46x36 = rnx46x35 || v32c;
wire onx46x36 = onx46x35 || ( rnx46x35 && v32c);
wire [16:0] v32d = 17'b11100110100101101;
wire v32e = v32d == v1c1;
wire v32f = v66 == v2d7;
wire v330 = v32e & v32f & v2c0 & v157 & v2ed;
wire v331 = v1ab == Advice_26;
wire v332 = Advice_19 == Advice_15;
wire v333 = v2d2 & v31 & v33 & v330 & v2d0 & v2b9 & v331 & v2cb & v2db & v2dd & v70 & v89 & v332 & v2f0 & v2ce;
wire rnx46x37 = rnx46x36 || v333;
wire onx46x37 = onx46x36 || ( rnx46x36 && v333);
wire v334 = v212 == Advice_14;
wire [15:0] v335 = 16'b0010011010010110;
wire v336 = v335 == vb7;
wire v337 = v336 & v218 & v326 & v9e & v2ed;
wire v339 = v212 == Advice_31;
wire [31:0] v33a = v203 + v10f;
wire [31:0] v33b = v33a + vab;
wire [31:0] v33c = v33b + vae;
wire v33d = v33c == Advice_26;
wire [2:0] v33e = { Advice_31 , v2f };
wire v33f = v33e == Advice_22;
wire v340 = v2b7 & v2a1 & v2b9 & v334 & v337 & v31 & v2cb & v339 & v70 & v33d & v33 & v89 & v173 & v33f & v2ce;
wire rnx46x38 = rnx46x37 || v340;
wire onx46x38 = onx46x37 || ( rnx46x37 && v340);
wire [2:0] v341 = instruction_bits[13: 11];
wire [2:0] v342 = { v341 };
wire v343 = v342 == Advice_6;
wire [31:0] v344 = v147 + vab;
wire [31:0] v345 = v344 + v14a;
wire v346 = v345 == Advice_26;
wire [10:0] v347 = 11'b10010110001;
wire [10:0] v348 = instruction_bits[10: 0];
wire v349 = v347 == v348;
wire [9:0] v34a = 10'b0010100101;
wire [9:0] v34b = instruction_bits[23: 14];
wire v34c = v34a == v34b;
wire v34d = v349 & v34c & v301 & v2ed;
wire v34e = v2f9 & v31 & v2b9 & v33 & v343 & v346 & v70 & v34d & v2f6 & v89 & v2ce;
wire rnx46x39 = rnx46x38 || v34e;
wire onx46x39 = onx46x38 || ( rnx46x38 && v34e);
wire [31:0] v34f = 32'b10010000000000000000000000000000;
wire [31:0] v350 = In_register_EIP + v34f;
wire v351 = v350 == Out_register_EIP;
wire v352 = v2aa & v2ab & v2ac & v2ad & v2ae & v2af & v2b0 & v2b1 & v351 & v50 & v51 & v52 & v53 & v54 & v55 & v56 & v2b4 & v5a & v2b5 & v5c & v5d & v5e;
wire v353 = v2a8 & v352;
wire [31:0] v354 = instruction_bits[71: 40];
wire v356 = v354 == Advice_24;
wire [31:0] v357 = v10f << v79;
wire [31:0] v358 = v75 + v357;
wire [31:0] v359 = v358 + v7e;
wire v35a = v359 == Advice_26;
wire v35c = instruction_bits[27: 27];
wire v35b = instruction_bits[29: 29];
wire [1:0] v35d = { v35c , v35b };
wire v35e = v35d == Advice_13;
wire v35f = instruction_bits[28: 28];
wire v360 = v66 == v35f;
wire [47:0] v361 = 48'b000000000000000000000000000000000000000000000000;
wire [47:0] v362 = instruction_bits[119: 72];
wire v363 = v361 == v362;
wire v364 = v2bf & v326 & v360 & v363 & v2ed;
wire v365 = Advice_13 == Advice_12;
wire v366 = v353 & v356 & v31 & v2bd & v2b9 & v35a & v2bc & v33 & v35e & v364 & v70 & v2cb & v89 & v145 & v365 & v2cd & v2ce;
wire rnx46x40 = rnx46x39 || v366;
wire onx46x40 = onx46x39 || ( rnx46x39 && v366);
wire [31:0] v367 = v204 + vab;
wire [31:0] v368 = v367 + va9;
wire v369 = v368 == Advice_26;
wire v36a = v68 & v2c1;
wire v36b = v36a ^ v66;
wire v36c = Advice_27 == v67;
wire v36d = v36c & v2c4;
wire v36e = v36d ^ v66;
wire v36f = v66 & v36b & v66 & v36e;
wire v370 = v336 & v2c0 & v157 & v36f;
wire v371 = Advice_27 == Advice_22;
wire v372 = v2d2 & v369 & v33 & v2b9 & v2d0 & v324 & v31 & v370 & v2cb & v89 & v328 & v70 & v145 & v371 & v2ce;
wire rnx46x41 = rnx46x40 || v372;
wire onx46x41 = onx46x40 || ( rnx46x40 && v372);
wire v373 = v292 == Advice_26;
wire [15:0] v374 = 16'b0110010010010110;
wire v375 = v374 == vb7;
wire v376 = v36c;
wire v377 = v376 ^ v66;
wire v378 = v66 & v6a & v66 & v377;
wire v379 = v375 & v310 & v301 & v378;
wire v37a = Advice_27 == Advice_8;
wire v37b = v2f9 & v31 & v33 & v2b9 & v2f6 & v324 & v89 & v328 & v373 & v379 & v2cb & v70 & v145 & v37a & v2ce;
wire rnx46x42 = rnx46x41 || v37b;
wire onx46x42 = onx46x41 || ( rnx46x41 && v37b);
wire [31:0] v37c = v31f + v1e9;
wire [15:0] v37d = v37c[15:0];
wire [31:0] v37e = { 16'b0000000000000000, v37d };
wire v37f = v37e == Advice_26;
wire v380 = v2d6 & v310 & v363 & v2ed;
wire v381 = v353 & v356 & v31 & v33 & vb4 & v2b9 & v324 & v37f & v2cb & v380 & v70 & v328 & v89 & v329 & v32a & v32b & v2ce;
wire rnx46x43 = rnx46x42 || v381;
wire onx46x43 = onx46x42 || ( rnx46x42 && v381);
wire v382 = ve5 == Advice_7;
wire [4:0] v383 = instruction_bits[18: 14];
wire v384 = vb9 == v383;
wire v385 = v349 & v384 & v301 & v314;
wire v386 = v14c == Advice_26;
wire v387 = Advice_7 == Advice_4;
wire v388 = v2f6 & v2f9 & v33 & v382 & v2b9 & v385 & v343 & v70 & v386 & v31 & v89 & v387 & v2ce;
wire rnx46x44 = rnx46x43 || v388;
wire onx46x44 = onx46x43 || ( rnx46x43 && v388);
wire [1:0] v389 = instruction_bits[15: 14];
wire v38a = v325 == v389;
wire v38b = v66 & v36b & v66 & v66;
wire v38c = v349 & v38a & vd1 & v9e & v38b;
wire v38d = vb0 == Advice_26;
wire v38e = Advice_27 == Advice_9;
wire v38f = v2b7 & v2a1 & v33 & v2b9 & v38c & v328 & v70 & v324 & v31 & v343 & v38d & v89 & v145 & v38e & v2ce;
wire rnx46x45 = rnx46x44 || v38f;
wire onx46x45 = onx46x44 || ( rnx46x44 && v38f);
wire v390 = vcc == Advice_26;
wire v391 = v1f7 == v389;
wire v392 = v66 & v36b & v66 & v2c6;
wire v393 = v349 & v391 & vd1 & v157 & v392;
wire v394 = v89 & v2d0 & v2d2 & v33 & v390 & v2b9 & v328 & v31 & v324 & v70 & v343 & v393 & v145 & v38e & v2ce;
wire rnx46x46 = rnx46x45 || v394;
wire onx46x46 = onx46x45 || ( rnx46x45 && v394);
wire v395 = v15a == Advice_26;
wire v396 = v2ea == v389;
wire v397 = v349 & v396 & vd1 & v301 & v38b;
wire v398 = v2f9 & v2f6 & v31 & v395 & v33 & v324 & v328 & v2b9 & v89 & v343 & v397 & v70 & v145 & v38e & v2ce;
wire rnx46x47 = rnx46x46 || v398;
wire onx46x47 = onx46x46 || ( rnx46x46 && v398);
wire [31:0] v399 = ve1 + v14a;
wire v39a = v399 == Advice_26;
wire v39b = v66 & v36b & v161 & v66;
wire v39c = v349 & v396 & v301 & v39b;
wire v39d = v39a & v2f9 & v33 & v2b9 & v324 & v31 & v382 & v2f6 & v328 & v39c & v343 & v70 & v89 & v145 & v2cc & v38e & v2ce;
wire rnx46x48 = rnx46x47 || v39d;
wire onx46x48 = onx46x47 || ( rnx46x47 && v39d);
wire v39e = ve2 == Advice_26;
wire v39f = v349 & v38a & v9e & v39b;
wire v3a0 = v2b7 & v39e & v2b9 & v33 & v382 & v328 & v2a1 & v39f & v324 & v343 & v70 & v31 & v89 & v145 & v2cc & v38e & v2ce;
wire rnx46x49 = rnx46x48 || v3a0;
wire onx46x49 = onx46x48 || ( rnx46x48 && v3a0);
wire v3a1 = v66 & v36b & v161 & v2c6;
wire v3a2 = v349 & v391 & v157 & v3a1;
wire [31:0] v3a3 = ve1 + va9;
wire v3a4 = v3a3 == Advice_26;
wire v3a5 = v2d2 & v2d0 & v3a2 & v3a4 & v89 & v33 & v31 & v70 & v2b9 & v324 & v328 & v343 & v382 & v145 & v2cc & v38e & v2ce;
wire rnx46x50 = rnx46x49 || v3a5;
wire onx46x50 = onx46x49 || ( rnx46x49 && v3a5);
wire [31:0] v3a6 = vac + v113;
wire v3a7 = v3a6 == Advice_26;
wire v3a8 = vef == Advice_27;
wire v3a9 = vef == Advice_2;
wire [7:0] v3aa = 8'b10010110;
wire v3ab = v3aa == vf3;
wire v3ac = v3ab & v38a & v157 & v378;
wire v3ad = v3a7 & v33 & v2b9 & v31 & v2d2 & v3a8 & v343 & v2d0 & v70 & v3a9 & v3ac & v89 & v145 & v38e & v2ce;
wire rnx46x51 = rnx46x50 || v3ad;
wire onx46x51 = onx46x50 || ( rnx46x50 && v3ad);
wire [31:0] v3ae = v344 + v17d;
wire v3af = v3ae == Advice_26;
wire [31:0] v3b0 = instruction_bits[79: 48];
wire v3b2 = v3b0 == Advice_24;
wire [10:0] v3b3 = 11'b10010110101;
wire v3b4 = v3b3 == v348;
wire [39:0] v3b5 = 40'b0000000000000000000000000000000000000000;
wire [39:0] v3b6 = instruction_bits[119: 80];
wire v3b7 = v3b5 == v3b6;
wire v3b8 = v3b4 & v391 & v3b7 & v2ed;
wire [31:0] v3b9 = 32'b01010000000000000000000000000000;
wire [31:0] v3ba = In_register_EIP + v3b9;
wire v3bb = v3ba == Out_register_EIP;
wire v3bc = v2aa & v2ab & v2ac & v2ad & v2ae & v2af & v2b0 & v2b1 & v3bb & v50 & v51 & v52 & v53 & v54 & v55 & v56 & v2b4 & v5a & v2b5 & v5c & v5d & v5e;
wire v3bd = v2a8 & v3bc;
wire v3be = v3af & v3b2 & v33 & v2b9 & v343 & v31 & v3b8 & v70 & v3bd & v89 & v2ce;
wire rnx46x52 = rnx46x51 || v3be;
wire onx46x52 = onx46x51 || ( rnx46x51 && v3be);
wire v3bf = v17d == Advice_24;
wire v3c0 = v2aa & v2ab & v2ac & v2ad & v2ae & v2af & v2b0 & v2b1 & v183 & v50 & v51 & v52 & v53 & v54 & v55 & v56 & v2b4 & v5a & v2b5 & v5c & v5d & v5e;
wire v3c1 = v2a8 & v3c0;
wire v3c2 = v3ab & v391 & v18a & v36f;
wire v3c3 = v3bf & v2b9 & v3a8 & v3c1 & v3a9 & v390 & v33 & v343 & v70 & v31 & v3c2 & v89 & v145 & v38e & v2ce;
wire rnx46x53 = rnx46x52 || v3c3;
wire onx46x53 = onx46x52 || ( rnx46x52 && v3c3);
wire [31:0] v3c4 = v111 + v17d;
wire v3c5 = v3c4 == Advice_26;
wire v3c6 = v109 == Advice_31;
wire v3c7 = v3ab & v102 & v396 & v3b7 & v2ed;
wire v3c8 = v109 == Advice_14;
wire v3c9 = Advice_31 == Advice_11;
wire v3ca = v3bd & v3c5 & v3c6 & v2b9 & v31 & v33 & v70 & v3c7 & v3c8 & v89 & v343 & v3b2 & v173 & v3c9 & v2ce;
wire rnx46x54 = rnx46x53 || v3ca;
wire onx46x54 = onx46x53 || ( rnx46x53 && v3ca);
wire v3cb =  v254 == memory_0[15: 12] && Advice_26 == memory_0[47: 16] && In_timestamp == memory_0[143: 80] && 4'd0 == memory_0[11: 8] && 1'b1 == memory_0[0: 0] && 6'b000000 == memory_0[7: 2] && 1'b0 == memory_0[1: 1];
wire [15:0] v3d0 = v77[31: 16];
wire [31:0] v3cc = Advice_24 << v248;
wire [31:0] v3cd = v3cc >>> v248;
wire [31:0] v3ce = v3cd * v23f;
wire [15:0] v3cf = v3ce[15:0];
wire [31:0] v3d1 = { v3d0 , v3cf };
wire v3d2 = v3d1 == v2a7;
wire [31:0] v3d3 = v3ce + v24e;
wire v3d4 = v3d3 < v23c;
wire v3d5 = v3d4 == Out_register_CF;
wire v3d6 = v3d4 == Out_register_OF;
wire v3d7 = v2aa & v2ab & v2ac & v2ad & v2ae & v2af & v2b0 & v2b1 & v183 & v50 & v51 & v52 & v53 & v54 & v55 & v56 & v3d5 & v5a & v3d6 & v5c & v5d & v5e;
wire v3d8 = v3d2 & v3d7;
wire [15:0] v3d9 = instruction_bits[47: 32];
wire [15:0] pad_986 = (v3d9[15:15] == 1'b1) ?16'b1111111111111111 : 16'b0000000000000000;
wire [31:0] v3da = { pad_986, v3d9 };
wire v3dc = v3da == Advice_24;
wire [18:0] v3dd = 19'b0110011010010110001;
wire v3de = v3dd == v153;
wire [4:0] v3df = instruction_bits[31: 27];
wire v3e0 = v103 == v3df;
wire v3e1 = v66 & v2c3 & v66 & v2c6;
wire v3e2 = v3de & v2c0 & v3e0 & v18a & v3e1;
wire v3e3 = Advice_6 == Advice_5;
wire v3e4 = v390 & v31 & v33 & v3cb & v2bd & v2bc & v3d8 & v2cb & v70 & v89 & v3dc & v3e2 & v145 & v38e & v2ce & v3e3;
wire rnx46x55 = rnx46x54 || v3e4;
wire onx46x55 = onx46x54 || ( rnx46x54 && v3e4);
wire [31:0] v3e6 = ( Advice_32 == 3'd0) ? In_register_EAX :
	( Advice_32 == 3'd1) ? In_register_ECX :
	( Advice_32 == 3'd2) ? In_register_EDX :
	( Advice_32 == 3'd3) ? In_register_EBX :
	( Advice_32 == 3'd4) ? In_register_ESP :
	( Advice_32 == 3'd5) ? In_register_EBP :
	( Advice_32 == 3'd6) ? In_register_ESI : In_register_EDI;
wire [15:0] v3e7 = v3e6[31: 16];
wire [31:0] v3e8 = { v3e7 , v3cf };
wire v3e9 = v3e8 == v2a7;
wire v3ea = v2aa & v2ab & v2ac & v2ad & v2ae & v2af & v2b0 & v2b1 & v150 & v50 & v51 & v52 & v53 & v54 & v55 & v56 & v3d5 & v5a & v3d6 & v5c & v5d & v5e;
wire v3eb = v3e9 & v3ea;
wire [15:0] v3ec = instruction_bits[55: 40];
wire [15:0] pad_1005 = (v3ec[15:15] == 1'b1) ?16'b1111111111111111 : 16'b0000000000000000;
wire [31:0] v3ed = { pad_1005, v3ec };
wire v3ef = v3ed == Advice_24;
wire v3f0 = v3de & v326 & v157 & v39b;
wire [31:0] v3f1 = va8 + v7b;
wire [31:0] v3f2 = v3f1 + v7e;
wire v3f3 = v3f2 == Advice_26;
wire v3f4 = Advice_6 == Advice_32;
wire v3f5 = v3eb & v3ef & v3cb & v31 & v33 & v2ba & v70 & v3f0 & v2bd & v2bc & v2cb & v3f3 & v89 & v145 & v2cc & v38e & v2ce & v3f4;
wire rnx46x56 = rnx46x55 || v3f5;
wire onx46x56 = onx46x55 || ( rnx46x55 && v3f5);
wire [15:0] v3f6 = 16'b0110011010010110;
wire v3f7 = v3f6 == vb7;
wire v3f8 = v66 & v36b & v66 & v377;
wire v3f9 = v3f7 & v326 & v18a & v3f8;
wire v3fa = v3d8 & v3dc & v89 & v38d & v3cb & v328 & v31 & v2cb & v33 & v70 & v324 & v3f9 & v145 & v38e & v2ce & v3e3;
wire rnx46x57 = rnx46x56 || v3fa;
wire onx46x57 = onx46x56 || ( rnx46x56 && v3fa);
wire [15:0] v3fb = v74[31: 16];
wire [31:0] v3fc = { v3fb , v3cf };
wire v3fd = v3fc == v2a7;
wire v3fe = v2aa & v2ab & v2ac & v2ad & v2ae & v2af & v2b0 & v2b1 & v4f & v50 & v51 & v52 & v53 & v54 & v55 & v56 & v3d5 & v5a & v3d6 & v5c & v5d & v5e;
wire v3ff = v3fd & v3fe;
wire v400 = v1e9 == Advice_24;
wire v401 = v20f == Advice_26;
wire v402 = v3f7 & v218 & v2c0 & v65 & v2ed;
wire v403 = v3ff & v400 & v31 & v401 & v3cb & v339 & v70 & v334 & v2cb & v402 & v33 & v89 & v173 & v3c9 & v2ce & v8a;
wire rnx46x58 = rnx46x57 || v403;
wire onx46x58 = onx46x57 || ( rnx46x57 && v403);
wire [15:0] v404 = instruction_bits[79: 64];
wire [15:0] pad_1029 = (v404[15:15] == 1'b1) ?16'b1111111111111111 : 16'b0000000000000000;
wire [31:0] v405 = { pad_1029, v404 };
wire v407 = v405 == Advice_24;
wire [31:0] v408 = v3f1 + v96;
wire v409 = v408 == Advice_26;
wire v40a = v3de & v310 & v3b7 & v39b;
wire v40b = v2aa & v2ab & v2ac & v2ad & v2ae & v2af & v2b0 & v2b1 & v3bb & v50 & v51 & v52 & v53 & v54 & v55 & v56 & v3d5 & v5a & v3d6 & v5c & v5d & v5e;
wire v40c = v3e9 & v40b;
wire v40d = v407 & v89 & v31 & v2bc & v409 & v33 & v2bd & v40a & v70 & v40c & v2cb & v3cb & v2ba & v145 & v2cc & v38e & v2ce & v3f4;
wire rnx46x59 = rnx46x58 || v40d;
wire onx46x59 = onx46x58 || ( rnx46x58 && v40d);
wire v40e = v3f7 & v310 & v363 & v378;
wire v40f = v2aa & v2ab & v2ac & v2ad & v2ae & v2af & v2b0 & v2b1 & v351 & v50 & v51 & v52 & v53 & v54 & v55 & v56 & v3d5 & v5a & v3d6 & v5c & v5d & v5e;
wire v410 = v3d2 & v40f;
wire [15:0] v411 = instruction_bits[71: 56];
wire [15:0] pad_1042 = (v411[15:15] == 1'b1) ?16'b1111111111111111 : 16'b0000000000000000;
wire [31:0] v412 = { pad_1042, v411 };
wire v414 = v412 == Advice_24;
wire v415 = v31 & v395 & v33 & v324 & v40e & v328 & v410 & v414 & v70 & v2cb & v3cb & v89 & v145 & v38e & v2ce & v3e3;
wire rnx46x60 = rnx46x59 || v415;
wire onx46x60 = onx46x59 || ( rnx46x59 && v415);
wire v416 = v7e == Advice_24;
wire [31:0] v417 = v93 + v10f;
wire [31:0] v418 = v417 + v11c;
wire [31:0] v419 = v418 + va9;
wire v41a = v419 == Advice_26;
wire [18:0] v41b = 19'b0110010011010110001;
wire v41c = v41b == v153;
wire v41d = v41c & v2c0 & v141 & v65 & v314;
wire v41e = v2aa & v2ab & v2ac & v2ad & v2ae & v2af & v2b0 & v2b1 & v4f & v50 & v51 & v52 & v53 & v54 & v55 & v56 & v2b4 & v5a & v2b5 & v5c & v5d & v5e;
wire v41f = v2a8 & v41e;
wire v420 = v13b == Advice_31;
wire v421 = v13b == Advice_14;
wire v422 = v33e == Advice_8;
wire v423 = v416 & v2cb & v41a & v31 & v70 & v2b9 & v41d & v2ba & v41f & v33 & v89 & v420 & v421 & v173 & v387 & v422 & v2ce;
wire rnx46x61 = rnx46x60 || v423;
wire onx46x61 = onx46x60 || ( rnx46x60 && v423);
wire v424 = v399 == Advice_1;
wire [15:0] v425 = 16'b0110111100110101;
wire v426 = v425 == vb7;
wire v427 = v426 & v157 & ve7;
wire v428 = v424 & v28c & v31 & v144 & v33 & v427 & v89 & ve6 & vb5 & vb4 & v70 & v8a & v8b & vc6;
wire rnx46x62 = rnx46x61 || v428;
wire onx46x62 = onx46x61 || ( rnx46x61 && v428);
wire v429 = v2aa & v2ab & v2ac & v2ad & v2ae & v2af & v2b0 & v2b1 & va4 & v50 & v51 & v52 & v53 & v54 & v55 & v56 & v2b4 & v5a & v2b5 & v5c & v5d & v5e;
wire v42a = v2a8 & v429;
wire [31:0] v42b = v1e7 + va9;
wire [15:0] v42c = v42b[15:0];
wire [31:0] v42d = { 16'b0000000000000000, v42c };
wire v42e = v42d == Advice_26;
wire [15:0] v42f = 16'b1110011011010110;
wire v430 = v42f == vb7;
wire v431 = Advice_19;
wire v432 = v431 ^ v66;
wire v433 = v66 & v432 & v66 & v66;
wire v434 = v430 & v2d8 & v2c0 & vbe & v433;
wire v435 = vae == Advice_24;
wire [2:0] v436 = { Advice_19 , v1f7 };
wire v437 = v436 == Advice_20;
wire v438 = v42a & v42e & v434 & v33 & v31 & v2b9 & v2dd & v435 & v2d4 & v2cb & v2db & v70 & v89 & v437 & v2df & v2e1 & v2ce;
wire rnx46x63 = rnx46x62 || v438;
wire onx46x63 = onx46x62 || ( rnx46x62 && v438);
wire [31:0] v439 = v1e7 + vae;
wire [15:0] v43a = v439[15:0];
wire [31:0] v43b = { 16'b0000000000000000, v43a };
wire v43c = v43b == Advice_26;
wire v43d = v430 & v2d8 & v326 & v65 & v433;
wire v43e = v41f & v416 & v2dd & v43c & v31 & v2cb & v33 & v89 & v2d4 & v2b9 & v43d & v70 & v2db & v437 & v2df & v2e1 & v2ce;
wire rnx46x64 = rnx46x63 || v43e;
wire onx46x64 = onx46x63 || ( rnx46x63 && v43e);
wire [16:0] v43f = 17'b11100110110101101;
wire v440 = v43f == v1c1;
wire v441 = v440 & v32f & v2c0 & vbe & v2ed;
wire v442 = v42a & v89 & v435 & v2dd & v2cb & v2b9 & v441 & v31 & v331 & v70 & v2db & v33 & v332 & v2f0 & v2ce;
wire rnx46x65 = rnx46x64 || v442;
wire onx46x65 = onx46x64 || ( rnx46x64 && v442);
wire [31:0] v443 = v205 + v7e;
wire v444 = v443 == Advice_26;
wire [18:0] v445 = 19'b0010011011010110001;
wire v446 = v445 == v153;
wire v447 = v446 & v326 & v18a & v314;
wire [7:0] v448 = instruction_bits[47: 40];
wire [7:0] pad_1097 = (v448[7:7] == 1'b1) ?24'b111111111111111111111111 : 24'b000000000000000000000000;
wire [31:0] v449 = { pad_1097, v448 };
wire v44b = v449 == Advice_24;
wire v44c = v3c1 & v31 & v2b9 & v33 & v2bd & v444 & v89 & v447 & v70 & v2bc & v2ba & v44b & v2cb & v145 & v2cc & v371 & v2ce;
wire rnx46x66 = rnx46x65 || v44c;
wire onx46x66 = onx46x65 || ( rnx46x65 && v44c);
wire [31:0] v44d = v291 + vae;
wire v44e = v44d == Advice_26;
wire [15:0] v44f = 16'b0110010011010110;
wire v450 = v44f == vb7;
wire v451 = v450 & v326 & v65 & v378;
wire v452 = v41f & v70 & v324 & v44e & v31 & v416 & v2b9 & v328 & v89 & v451 & v33 & v2cb & v145 & v37a & v2ce;
wire rnx46x67 = rnx46x66 || v452;
wire onx46x67 = onx46x66 || ( rnx46x66 && v452);
wire v453 = v450 & v218 & v2c0 & vbe & v2ed;
wire [31:0] v454 = v417 + vab;
wire [31:0] v455 = v454 + va9;
wire v456 = v455 == Advice_26;
wire v457 = v435 & v453 & v31 & v42a & v33 & v2cb & v334 & v2b9 & v70 & v456 & v339 & v89 & v173 & v422 & v2ce;
wire rnx46x68 = rnx46x67 || v457;
wire onx46x68 = onx46x67 || ( rnx46x67 && v457);
wire [31:0] v458 = In_register_FSBASE + va9;
wire [31:0] v459 = v458 + vab;
wire [31:0] v45a = v459 + v14a;
wire v45b = v45a == Advice_26;
wire [18:0] v45c = 19'b0010011011010110101;
wire v45d = v45c == v153;
wire v45e = v45d & v2c0 & v9e & v2ed;
wire [7:0] v45f = instruction_bits[63: 56];
wire [7:0] pad_1120 = (v45f[7:7] == 1'b1) ?24'b111111111111111111111111 : 24'b000000000000000000000000;
wire [31:0] v460 = { pad_1120, v45f };
wire v462 = v460 == Advice_24;
wire v463 = v2b7 & v45b & v31 & v2b9 & v2cb & v45e & v70 & v462 & v33 & v89 & v2ce;
wire rnx46x69 = rnx46x68 || v463;
wire onx46x69 = onx46x68 || ( rnx46x68 && v463);
wire [10:0] v464 = 11'b11010110001;
wire v465 = v464 == v348;
wire [9:0] v466 = 10'b0010100111;
wire v467 = v466 == v34b;
wire v468 = v465 & v467 & v9e & v2ed;
wire v469 = v462 & v346 & v33 & v343 & v2b7 & v468 & v70 & v2b9 & v31 & v89 & v2ce;
wire rnx46x70 = rnx46x69 || v469;
wire onx46x70 = onx46x69 || ( rnx46x69 && v469);
wire [7:0] v46a = instruction_bits[71: 64];
wire [7:0] pad_1131 = (v46a[7:7] == 1'b1) ?24'b111111111111111111111111 : 24'b000000000000000000000000;
wire [31:0] v46b = { pad_1131, v46a };
wire v46d = v46b == Advice_24;
wire v46e = v98 == Advice_26;
wire v46f = v41c & v310 & v363 & v314;
wire v470 = v353 & v46d & v70 & v2b9 & v2bc & v2bd & v2cb & v33 & v89 & v46e & v2ba & v46f & v31 & v145 & v2cc & v37a & v2ce;
wire rnx46x71 = rnx46x70 || v470;
wire onx46x71 = onx46x70 || ( rnx46x70 && v470);
wire v471 = v1ed == Advice_26;
wire v472 = v430 & v2d8 & v310 & v18a & v433;
wire v473 = v3c1 & v44b & v31 & v33 & v471 & v2b9 & v2dd & v70 & v2db & v2d4 & v2cb & v472 & v89 & v437 & v2df & v2e1 & v2ce;
wire rnx46x72 = rnx46x71 || v473;
wire onx46x72 = onx46x71 || ( rnx46x71 && v473);
wire v474 = v450 & v310 & v9e & v378;
wire v475 = v2b7 & v462 & v89 & v31 & v373 & v328 & v324 & v70 & v2cb & v33 & v2b9 & v474 & v145 & v37a & v2ce;
wire rnx46x73 = rnx46x72 || v475;
wire onx46x73 = onx46x72 || ( rnx46x72 && v475);
wire v476 = v465 & v38a & vd1 & v65 & v38b;
wire v477 = v41f & v343 & v38d & v31 & v33 & v324 & v476 & v328 & v416 & v2b9 & v70 & v89 & v145 & v38e & v2ce;
wire rnx46x74 = rnx46x73 || v477;
wire onx46x74 = onx46x73 || ( rnx46x73 && v477);
wire v478 = v465 & v391 & vd1 & vbe & v392;
wire v479 = v390 & v42a & v33 & v31 & v2b9 & v435 & v324 & v328 & v343 & v478 & v70 & v89 & v145 & v38e & v2ce;
wire rnx46x75 = rnx46x74 || v479;
wire onx46x75 = onx46x74 || ( rnx46x74 && v479);
wire v47a = v465 & v396 & vd1 & v9e & v38b;
wire v47b = v462 & v70 & v31 & v2b9 & v343 & v2b7 & v328 & v395 & v89 & v33 & v47a & v324 & v145 & v38e & v2ce;
wire rnx46x76 = rnx46x75 || v47b;
wire onx46x76 = onx46x75 || ( rnx46x75 && v47b);
wire v47c = v16c == Advice_13;
wire [31:0] v47d = v147 + v16f;
wire [31:0] v47e = v47d + v14a;
wire v47f = v47e == Advice_26;
wire v480 = v465 & v384 & v168 & v9e & v2ed;
wire v481 = v2b7 & v462 & v33 & v2b9 & v47c & v343 & v47f & v31 & v480 & v70 & v89 & v365 & v2ce;
wire rnx46x77 = rnx46x76 || v481;
wire onx46x77 = onx46x76 || ( rnx46x76 && v481);
wire v482 = Advice_2 == v21d;
wire v483 = Advice_2 == v21f;
wire v484 = Advice_2 == v221;
wire v485 = Advice_2 == v223;
wire v486 = Advice_2 == v225;
wire v487 = Advice_2 == v227;
wire v488 = v482 & v483 & v484 & v485 & v486 & v487;
wire v489 = v488 ^ v66;
wire v48a = v66 & v489 & v161 & v66;
wire v48b = v465 & v38a & v65 & v48a;
wire v48c = v41f & v39e & v31 & v2b9 & v382 & v89 & v70 & v328 & v48b & v33 & v324 & v416 & v343 & v145 & v2cc & v38e & v2ce;
wire rnx46x78 = rnx46x77 || v48c;
wire onx46x78 = onx46x77 || ( rnx46x77 && v48c);
wire v48d = v465 & v396 & v9e & v48a;
wire v48e = v2b7 & v39a & v89 & v31 & v2b9 & v324 & v33 & v328 & v343 & v462 & v382 & v48d & v70 & v145 & v2cc & v38e & v2ce;
wire rnx46x79 = rnx46x78 || v48e;
wire onx46x79 = onx46x78 || ( rnx46x78 && v48e);
wire v48f = v465 & v391 & vbe & v3a1;
wire v490 = v435 & v31 & v42a & v2b9 & v48f & v33 & v324 & v3a4 & v382 & v328 & v343 & v70 & v89 & v145 & v2cc & v38e & v2ce;
wire rnx46x80 = rnx46x79 || v490;
wire onx46x80 = onx46x79 || ( rnx46x79 && v490);
wire [7:0] v491 = instruction_bits[55: 48];
wire [7:0] pad_1170 = (v491[7:7] == 1'b1) ?24'b111111111111111111111111 : 24'b000000000000000000000000;
wire [31:0] v492 = { pad_1170, v491 };
wire v494 = v492 == Advice_24;
wire [10:0] v495 = 11'b11010110101;
wire v496 = v495 == v348;
wire v497 = v496 & v391 & v157 & v2ed;
wire v498 = v2d2 & v3af & v31 & v2b9 & v494 & v33 & v70 & v497 & v343 & v89 & v2ce;
wire rnx46x81 = rnx46x80 || v498;
wire onx46x81 = onx46x80 || ( rnx46x80 && v498);
wire v499 = v17f == Advice_26;
wire [7:0] v49a = 8'b11010110;
wire v49b = v49a == vf3;
wire v49c = v49b & v396 & v157 & v3f8;
wire v49d = v2d2 & v499 & v33 & v49c & v2b9 & v494 & v89 & v3a9 & v3a8 & v31 & v343 & v70 & v145 & v38e & v2ce;
wire rnx46x82 = rnx46x81 || v49d;
wire onx46x82 = onx46x81 || ( rnx46x81 && v49d);
wire v49e = v49b & v38a & vbe & v378;
wire v49f = v42a & v3a7 & v31 & v2b9 & v3a8 & v343 & v49e & v435 & v70 & v3a9 & v33 & v89 & v145 & v38e & v2ce;
wire rnx46x83 = rnx46x82 || v49f;
wire onx46x83 = onx46x82 || ( rnx46x82 && v49f);
wire v4a0 = v2aa & v2ab & v2ac & v2ad & v2ae & v2af & v2b0 & v2b1 & vca & v50 & v51 & v52 & v53 & v54 & v55 & v56 & v2b4 & v5a & v2b5 & v5c & v5d & v5e;
wire v4a1 = v2a8 & v4a0;
wire v4a2 = v113 == Advice_24;
wire v4a3 = v49b & v391 & vd4 & v36f;
wire v4a4 = v4a1 & v4a2 & v31 & v33 & v343 & v2b9 & v3a8 & v89 & v390 & v3a9 & v4a3 & v70 & v145 & v38e & v2ce;
wire rnx46x84 = rnx46x83 || v4a4;
wire onx46x84 = onx46x83 || ( rnx46x83 && v4a4);
wire [31:0] pad_1189 = (Advice_26[31:31] == 1'b1) ?32'b11111111111111111111111111111111 : 32'b00000000000000000000000000000000;
wire [63:0] v4a5 = { pad_1189, Advice_26 };
wire [63:0] v4a6 = v2a2 * v4a5;
wire [31:0] v4a7 = v4a6[31:0];
wire [31:0] v4a8 = { v4a7 };
wire v4a9 = v4a8 == v2a7;
wire [63:0] v4aa = v4a6 + v1b5;
wire v4ab = v4aa < v1b7;
wire v4ac = v4ab == Out_register_CF;
wire v4ad = v4ab == Out_register_OF;
wire v4ae = v2aa & v2ab & v2ac & v2ad & v2ae & v2af & v2b0 & v2b1 & v90 & v50 & v51 & v52 & v53 & v54 & v55 & v56 & v4ac & v5a & v4ad & v5c & v5d & v5e;
wire v4af = v4a9 & v4ae;
wire v4b0 = v3a == Advice_6;
wire v4b1 = v74 == Advice_26;
wire [23:0] v4b2 = 24'b101001100010011010010110;
wire v4b3 = v4b2 == v61;
wire [1:0] v4b4 = 2'b11;
wire v4b5 = v4b4 == v78;
wire v4b6 = v66 & v66;
wire v4b7 = v4b3 & v4b5 & v9e & v4b6;
wire v4b8 = v31 & v4af & v33 & v2a1 & v2bd & v4b0 & v70 & v4b1 & v4b7 & v89 & v145 & v2ce;
wire rnx46x85 = rnx46x84 || v4b8;
wire onx46x85 = onx46x84 || ( rnx46x84 && v4b8);
wire v4b9 = v2aa & v2ab & v2ac & v2ad & v2ae & v2af & v2b0 & v2b1 & v150 & v50 & v51 & v52 & v53 & v54 & v55 & v56 & v4ac & v5a & v4ad & v5c & v5d & v5e;
wire v4ba = v4a9 & v4b9;
wire v4bb = v4b4 == vdd;
wire v4bc = v2d6 & v4bb & v157 & v4b6;
wire v4bd = v4ba & v2d0 & v33 & v328 & v70 & v2cb & v4b1 & v4bc & v31 & v89 & v145 & v2ce;
wire rnx46x86 = rnx46x85 || v4bd;
wire onx46x86 = onx46x85 || ( rnx46x85 && v4bd);
wire v4be = v2aa & v2ab & v2ac & v2ad & v2ae & v2af & v2b0 & v2b1 & v183 & v50 & v51 & v52 & v53 & v54 & v55 & v56 & v4ac & v5a & v4ad & v5c & v5d & v5e;
wire v4bf = v4a9 & v4be;
wire v4c0 = v4b4 == v389;
wire v4c1 = v3ab & v4c0 & v18a & v4b6;
wire v4c2 = v4bf & v3bf & v31 & v4b1 & v33 & v3a9 & v343 & v4c1 & v70 & v89 & v145 & v2ce;
wire rnx46x87 = rnx46x86 || v4c2;
wire onx46x87 = onx46x86 || ( rnx46x86 && v4c2);
wire [31:0] v4c3 = Advice_26 << v248;
wire [31:0] v4c4 = v4c3 >>> v248;
wire [31:0] v4c5 = v3cd * v4c4;
wire [15:0] v4c6 = v4c5[15:0];
wire [31:0] v4c7 = { v3d0 , v4c6 };
wire v4c8 = v4c7 == v2a7;
wire [31:0] v4c9 = v4c5 + v24e;
wire v4ca = v4c9 < v23c;
wire v4cb = v4ca == Out_register_CF;
wire v4cc = v4ca == Out_register_OF;
wire v4cd = v2aa & v2ab & v2ac & v2ad & v2ae & v2af & v2b0 & v2b1 & v183 & v50 & v51 & v52 & v53 & v54 & v55 & v56 & v4cb & v5a & v4cc & v5c & v5d & v5e;
wire v4ce = v4c8 & v4cd;
wire [31:0] v4cf = v74 & v1a5;
wire v4d0 = v4cf == Advice_26;
wire [23:0] v4d1 = 24'b011001000110011010010110;
wire v4d2 = v4d1 == v61;
wire v4d3 = v4d2 & v4b5 & v18a & v4b6;
wire v4d4 = v3dc & v31 & v33 & v2bd & v70 & v4ce & v4d0 & v4b0 & v4d3 & v89 & v145 & v2ce & v3e3;
wire rnx46x88 = rnx46x87 || v4d4;
wire onx46x88 = onx46x87 || ( rnx46x87 && v4d4);
wire v4d5 = v3f7 & v4bb & v65 & v4b6;
wire v4d6 = v2aa & v2ab & v2ac & v2ad & v2ae & v2af & v2b0 & v2b1 & v4f & v50 & v51 & v52 & v53 & v54 & v55 & v56 & v4cb & v5a & v4cc & v5c & v5d & v5e;
wire v4d7 = v4c8 & v4d6;
wire v4d8 = v4d0 & v31 & v33 & v4d5 & v328 & v2cb & v70 & v4d7 & v400 & v89 & v145 & v2ce & v3e3;
wire rnx46x89 = rnx46x88 || v4d8;
wire onx46x89 = onx46x88 || ( rnx46x88 && v4d8);
wire v4d9 = v2aa & v2ab & v2ac & v2ad & v2ae & v2af & v2b0 & v2b1 & v4f & v50 & v51 & v52 & v53 & v54 & v55 & v56 & v4ac & v5a & v4ad & v5c & v5d & v5e;
wire v4da = v4a9 & v4d9;
wire [23:0] v4db = 24'b101001101110011011010110;
wire v4dc = v4db == v61;
wire v4dd = v4dc & v4b5 & v65 & v4b6;
wire v4de = v4da & v416 & v4b1 & v31 & v33 & v89 & v4dd & v2bd & v4b0 & v70 & v145 & v2ce;
wire rnx46x90 = rnx46x89 || v4de;
wire onx46x90 = onx46x89 || ( rnx46x89 && v4de);
wire v4df = v2aa & v2ab & v2ac & v2ad & v2ae & v2af & v2b0 & v2b1 & va4 & v50 & v51 & v52 & v53 & v54 & v55 & v56 & v4ac & v5a & v4ad & v5c & v5d & v5e;
wire v4e0 = v4a9 & v4df;
wire v4e1 = v450 & v4bb & vbe & v4b6;
wire v4e2 = v4e0 & v435 & v4b1 & v31 & v33 & v2cb & v328 & v4e1 & v70 & v89 & v145 & v2ce;
wire rnx46x91 = rnx46x90 || v4e2;
wire onx46x91 = onx46x90 || ( rnx46x90 && v4e2);
wire v4e3 = v2aa & v2ab & v2ac & v2ad & v2ae & v2af & v2b0 & v2b1 & vca & v50 & v51 & v52 & v53 & v54 & v55 & v56 & v4ac & v5a & v4ad & v5c & v5d & v5e;
wire v4e4 = v4a9 & v4e3;
wire v4e5 = v49b & v4c0 & vd4 & v4b6;
wire v4e6 = v4a2 & v4e4 & v31 & v33 & v3a9 & v70 & v343 & v4e5 & v4b1 & v89 & v145 & v2ce;
wire rnx46x92 = rnx46x91 || v4e6;
wire onx46x92 = onx46x91 || ( rnx46x91 && v4e6);
wire [31:0] pad_1255 = (Advice_1[31:31] == 1'b1) ?32'b11111111111111111111111111111111 : 32'b00000000000000000000000000000000;
wire [63:0] v4e7 = { pad_1255, Advice_1 };
wire [63:0] v4e8 = v1ae * v4e7;
wire [31:0] v4e9 = v4e8[31:0];
wire v4ea = v4e9 == Out_register_EAX;
wire [63:0] v4eb = v4e8 >> v45;
wire [31:0] v4ec = v4eb[31:0];
wire v4ed = v4ec == Out_register_EDX;
wire [63:0] v4ee = v4e8 + v1b5;
wire v4ef = v4ee < v1b7;
wire v4f0 = v4ef == Out_register_CF;
wire v4f1 = v4ef == Out_register_OF;
wire v4f2 = v4ea & v43 & v44 & v4ed & v49 & v4a & v4b & v4c & vca & v50 & v51 & v52 & v53 & v54 & v55 & v56 & v4f0 & v5a & v4f1 & v5c & v5d & v5e;
wire [4:0] v4f3 = 5'b10111;
wire v4f4 = v4f3 == vba;
wire v4f5 = v1f0 & v4f4 & vd4 & v19c;
wire v4f6 = v4f2 & v199 & v31 & v33 & vb5 & v4f5 & v70 & v89 & v8a;
wire rnx46x93 = rnx46x92 || v4f6;
wire onx46x93 = onx46x92 || ( rnx46x92 && v4f6);
wire v4f7 = v4f3 == vf6;
wire v4f8 = vf4 & v4f7 & vfa & v19c;
wire v4f9 = v4ea & v43 & v44 & v4ed & v49 & v4a & v4b & v4c & vec & v50 & v51 & v52 & v53 & v54 & v55 & v56 & v4f0 & v5a & v4f1 & v5c & v5d & v5e;
wire v4fa = v33 & v4f8 & v4f9 & v70 & vf0 & v199 & v31 & v89 & v8a;
wire rnx46x94 = rnx46x93 || v4fa;
wire onx46x94 = onx46x93 || ( rnx46x93 && v4fa);
wire [31:0] v4fb = Advice_1 << v248;
wire [31:0] v4fc = v4fb >>> v248;
wire [31:0] v4fd = v4fc * v241;
wire [15:0] v4fe = v4fd[15:0];
wire [31:0] v4ff = { 16'b0000000000000000, v4fe };
wire [31:0] v500 = v23d | v4ff;
wire v501 = v500 == Out_register_EAX;
wire [31:0] v502 = v4fd >> v248;
wire [15:0] v503 = v502[15:0];
wire [31:0] v504 = { 16'b0000000000000000, v503 };
wire [31:0] v505 = v247 | v504;
wire v506 = v505 == Out_register_EDX;
wire [31:0] v507 = v4fd + v24e;
wire v508 = v507 < v23c;
wire v509 = v508 == Out_register_CF;
wire v50a = v508 == Out_register_OF;
wire v50b = v501 & v43 & v44 & v506 & v49 & v4a & v4b & v4c & va4 & v50 & v51 & v52 & v53 & v54 & v55 & v56 & v509 & v5a & v50a & v5c & v5d & v5e;
wire v50c = v4cf == Advice_1;
wire [23:0] v50d = 24'b011001100110011011101111;
wire v50e = v50d == v61;
wire v50f = v4f3 == v3df;
wire v510 = v50e & v50f & vbe & v19c;
wire v511 = v50b & v50c & v33 & v85 & v70 & v31 & v510 & v89 & v8a;
wire rnx46x95 = rnx46x94 || v511;
wire onx46x95 = onx46x94 || ( rnx46x94 && v511);
wire v512 = v3ae == Advice_1;
wire [15:0] v513 = 16'b0110111110100100;
wire v514 = v513 == vb7;
wire v515 = v514 & v18a & v105;
wire v516 = v184 & v512 & v31 & v144 & v70 & v515 & v33 & v89;
wire rnx46x96 = rnx46x95 || v516;
wire onx46x96 = onx46x95 || ( rnx46x95 && v516);
wire v517 = v345 == Advice_1;
wire v518 = v1b1 & v43 & v44 & v1b4 & v49 & v4a & v4b & v4c & v150 & v50 & v51 & v52 & v53 & v54 & v55 & v56 & v1b9 & v5a & v1ba & v5c & v5d & v5e;
wire [23:0] v519 = 24'b111011110011010010100110;
wire v51a = v519 == v61;
wire v51b = v51a & v157 & v105;
wire v51c = v517 & v518 & v31 & v33 & v51b & v38 & v70 & v89;
wire rnx46x97 = rnx46x96 || v51c;
wire onx46x97 = onx46x96 || ( rnx46x96 && v51c);
wire [15:0] v51d = 16'b1110111110110100;
wire v51e = v51d == vb7;
wire v51f = v51e & v18a & v105;
wire v520 = v512 & v33 & v51f & v31 & v70 & v38 & v237 & v89;
wire rnx46x98 = rnx46x97 || v520;
wire onx46x98 = onx46x97 || ( rnx46x97 && v520);
wire [31:0] v521 = v344 + v96;
wire v522 = v521 == Advice_1;
wire [31:0] v523 = 32'b01100110011001101110111110110100;
wire [31:0] v524 = instruction_bits[31: 0];
wire v525 = v523 == v524;
wire v526 = v525 & v9e & v105;
wire v527 = v246 & v43 & v44 & v24d & v49 & v4a & v4b & v4c & v90 & v50 & v51 & v52 & v53 & v54 & v55 & v56 & v251 & v5a & v252 & v5c & v5d & v5e;
wire v528 = v522 & v31 & v255 & v526 & v527 & v33 & v70 & v89;
wire rnx46x99 = rnx46x98 || v528;
wire onx46x99 = onx46x98 || ( rnx46x98 && v528);
wire v2e = (!onx46x99) && rnx46x99;
assign result = v2e;
assign dummy = 1'b0;
endmodule
