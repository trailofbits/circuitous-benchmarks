module circuit(
input [1726:0] current,
input [1726:0] next,

output [0:0] result,
output [0:0] dummy
);
wire Advice_1 = current[0: 0];
wire [31:0] Advice_10 = current[32: 1];
wire [2:0] Advice_11 = current[35: 33];
wire [2:0] Advice_12 = current[38: 36];
wire [2:0] Advice_13 = current[41: 39];
wire [2:0] Advice_14 = current[44: 42];
wire [1:0] Advice_15 = current[46: 45];
wire [1:0] Advice_16 = current[48: 47];
wire [2:0] Advice_17 = current[51: 49];
wire [2:0] Advice_18 = current[54: 52];
wire Advice_19 = current[55: 55];
wire [2:0] Advice_2 = current[58: 56];
wire Advice_20 = current[59: 59];
wire Advice_21 = current[60: 60];
wire [1:0] Advice_22 = current[62: 61];
wire [1:0] Advice_23 = current[64: 63];
wire [2:0] Advice_24 = current[67: 65];
wire [1:0] Advice_25 = current[69: 68];
wire Advice_26 = current[70: 70];
wire [2:0] Advice_27 = current[73: 71];
wire [2:0] Advice_28 = current[76: 74];
wire [2:0] Advice_29 = current[79: 77];
wire [2:0] Advice_3 = current[82: 80];
wire [2:0] Advice_30 = current[85: 83];
wire [2:0] Advice_31 = current[88: 86];
wire [1:0] Advice_32 = current[90: 89];
wire [31:0] Advice_4 = current[122: 91];
wire [31:0] Advice_5 = current[154: 123];
wire [2:0] Advice_6 = current[157: 155];
wire [2:0] Advice_7 = current[160: 158];
wire Advice_8 = current[161: 161];
wire Advice_9 = current[162: 162];
wire In_error_flag = current[163: 163];
wire In_register_AF = current[492: 492];
wire [31:0] In_register_CSBASE = current[525: 494];
wire [7:0] In_register_DF = current[533: 526];
wire [31:0] In_register_DSBASE = current[565: 534];
wire [31:0] In_register_EAX = current[597: 566];
wire [31:0] In_register_EBP = current[629: 598];
wire [31:0] In_register_EBX = current[661: 630];
wire [31:0] In_register_ECX = current[693: 662];
wire [31:0] In_register_EDI = current[725: 694];
wire [31:0] In_register_EDX = current[757: 726];
wire [31:0] In_register_EIP = current[789: 758];
wire [31:0] In_register_ESBASE = current[821: 790];
wire [31:0] In_register_ESI = current[853: 822];
wire [31:0] In_register_ESP = current[885: 854];
wire [31:0] In_register_FSBASE = current[917: 886];
wire [31:0] In_register_GSBASE = current[949: 918];
wire In_register_PF = current[951: 951];
wire In_register_SF = current[952: 952];
wire [31:0] In_register_SSBASE = current[984: 953];
wire In_register_ZF = current[985: 985];
wire [63:0] In_timestamp = current[1049: 986];
wire Out_error_flag = next[163: 163];
wire Out_register_AF = next[492: 492];
wire Out_register_CF = next[493: 493];
wire [31:0] Out_register_CSBASE = next[525: 494];
wire [7:0] Out_register_DF = next[533: 526];
wire [31:0] Out_register_DSBASE = next[565: 534];
wire [31:0] Out_register_EAX = next[597: 566];
wire [31:0] Out_register_EBP = next[629: 598];
wire [31:0] Out_register_EBX = next[661: 630];
wire [31:0] Out_register_ECX = next[693: 662];
wire [31:0] Out_register_EDI = next[725: 694];
wire [31:0] Out_register_EDX = next[757: 726];
wire [31:0] Out_register_EIP = next[789: 758];
wire [31:0] Out_register_ESBASE = next[821: 790];
wire [31:0] Out_register_ESI = next[853: 822];
wire [31:0] Out_register_ESP = next[885: 854];
wire [31:0] Out_register_FSBASE = next[917: 886];
wire [31:0] Out_register_GSBASE = next[949: 918];
wire Out_register_OF = next[950: 950];
wire Out_register_PF = next[951: 951];
wire Out_register_SF = next[952: 952];
wire [31:0] Out_register_SSBASE = next[984: 953];
wire Out_register_ZF = next[985: 985];
wire [63:0] Out_timestamp = next[1049: 986];
wire [119:0] instruction_bits = current[283: 164];
wire [207:0] memory_0 = current[491: 284];
wire [31:0] v4 = 32'b00000000000000001111111111111111;
wire [31:0] v5 = In_register_EAX & v4;
wire [15:0] v6 = 16'b1110011001101111;
wire [15:0] v8 = instruction_bits[15: 0];
wire v9 = v6 == v8;
wire [5:0] va = 6'b010110;
wire [5:0] vb = instruction_bits[23: 18];
wire vc = va == vb;
wire [87:0] vd = 88'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
wire [87:0] ve = instruction_bits[119: 32];
wire vf = vd == ve;
wire v11 = 1'b0;
wire v12 = Advice_1 == v11;
wire v13 = v12;
wire v14 = 1'b1;
wire v15 = v13 ^ v14;
wire v16 = v15 & v14 & v14;
wire v17 = v9 & vc & vf & v16;
wire v18 = v17;
wire [63:0] v19 = { v18 , v18 , v18 , v18 , v18 , v18 , v18 , v18 , v18 , v18 , v18 , v18 , v18 , v18 , v18 , v18 , v18 , v18 , v18 , v18 , v18 , v18 , v18 , v18 , v18 , v18 , v18 , v18 , v18 , v18 , v18 , v18 , v18 , v18 , v18 , v18 , v18 , v18 , v18 , v18 , v18 , v18 , v18 , v18 , v18 , v18 , v18 , v18 , v18 , v18 , v18 , v18 , v18 , v18 , v18 , v18 , v18 , v18 , v18 , v18 , v18 , v18 , v18 , v18 };
wire [31:0] v1b = memory_0[79: 48];
wire [7:0] v1c = v1b[7:0];
wire [7:0] pad_29 = (v1c[7:7] == 1'b1) ?8'b11111111 : 8'b00000000;
wire [15:0] v1d = { pad_29, v1c };
wire [15:0] pad_30 = (v1d[15:15] == 1'b1) ?48'b111111111111111111111111111111111111111111111111 : 48'b000000000000000000000000000000000000000000000000;
wire [63:0] v1e = { pad_30, v1d };
wire [63:0] v1f = v19 & v1e;
wire [15:0] v20 = 16'b0110111100100100;
wire v21 = v20 == v8;
wire v22 = instruction_bits[20: 20];
wire v23 = v14 == v22;
wire [95:0] v24 = 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
wire [95:0] v25 = instruction_bits[119: 24];
wire v26 = v24 == v25;
wire [2:0] v28 = 3'b101;
wire v29 = Advice_2 == v28;
wire v2a = v29;
wire v2b = v2a ^ v14;
wire v2c = v14 & v14 & v2b;
wire v2d = v21 & v23 & v26 & v2c;
wire v2e = v2d;
wire [63:0] v2f = { v2e , v2e , v2e , v2e , v2e , v2e , v2e , v2e , v2e , v2e , v2e , v2e , v2e , v2e , v2e , v2e , v2e , v2e , v2e , v2e , v2e , v2e , v2e , v2e , v2e , v2e , v2e , v2e , v2e , v2e , v2e , v2e , v2e , v2e , v2e , v2e , v2e , v2e , v2e , v2e , v2e , v2e , v2e , v2e , v2e , v2e , v2e , v2e , v2e , v2e , v2e , v2e , v2e , v2e , v2e , v2e , v2e , v2e , v2e , v2e , v2e , v2e , v2e , v2e };
wire [15:0] v30 = { 8'b00000000, v1c };
wire [15:0] pad_49 = (v30[15:15] == 1'b1) ?48'b111111111111111111111111111111111111111111111111 : 48'b000000000000000000000000000000000000000000000000;
wire [63:0] v31 = { pad_49, v30 };
wire [63:0] v32 = v2f & v31;
wire [15:0] v33 = 16'b0110111100100101;
wire v34 = v33 == v8;
wire [63:0] v35 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
wire [63:0] v36 = instruction_bits[119: 56];
wire v37 = v35 == v36;
wire v38 = v14 & v14 & v14;
wire v39 = v34 & v23 & v37 & v38;
wire v3a = v39;
wire [63:0] v3b = { v3a , v3a , v3a , v3a , v3a , v3a , v3a , v3a , v3a , v3a , v3a , v3a , v3a , v3a , v3a , v3a , v3a , v3a , v3a , v3a , v3a , v3a , v3a , v3a , v3a , v3a , v3a , v3a , v3a , v3a , v3a , v3a , v3a , v3a , v3a , v3a , v3a , v3a , v3a , v3a , v3a , v3a , v3a , v3a , v3a , v3a , v3a , v3a , v3a , v3a , v3a , v3a , v3a , v3a , v3a , v3a , v3a , v3a , v3a , v3a , v3a , v3a , v3a , v3a };
wire [63:0] v3c = v3b & v31;
wire [15:0] v3d = 16'b0110111110100100;
wire v3e = v3d == v8;
wire [71:0] v3f = 72'b000000000000000000000000000000000000000000000000000000000000000000000000;
wire [71:0] v40 = instruction_bits[119: 48];
wire v41 = v3f == v40;
wire v42 = v3e & v41 & v38;
wire v43 = v42;
wire [63:0] v44 = { v43 , v43 , v43 , v43 , v43 , v43 , v43 , v43 , v43 , v43 , v43 , v43 , v43 , v43 , v43 , v43 , v43 , v43 , v43 , v43 , v43 , v43 , v43 , v43 , v43 , v43 , v43 , v43 , v43 , v43 , v43 , v43 , v43 , v43 , v43 , v43 , v43 , v43 , v43 , v43 , v43 , v43 , v43 , v43 , v43 , v43 , v43 , v43 , v43 , v43 , v43 , v43 , v43 , v43 , v43 , v43 , v43 , v43 , v43 , v43 , v43 , v43 , v43 , v43 };
wire [63:0] v45 = v44 & v31;
wire [7:0] v46 = 8'b01101111;
wire [7:0] v47 = instruction_bits[7: 0];
wire v48 = v46 == v47;
wire [4:0] v49 = 5'b00101;
wire [4:0] v4a = instruction_bits[15: 11];
wire v4b = v49 == v4a;
wire [2:0] v4c = 3'b001;
wire v4d = Advice_2 == v4c;
wire v4e = v4d;
wire v4f = v4e ^ v14;
wire v50 = v14 & v14 & v4f;
wire v51 = v48 & v4b & v41 & v50;
wire v52 = v51;
wire [63:0] v53 = { v52 , v52 , v52 , v52 , v52 , v52 , v52 , v52 , v52 , v52 , v52 , v52 , v52 , v52 , v52 , v52 , v52 , v52 , v52 , v52 , v52 , v52 , v52 , v52 , v52 , v52 , v52 , v52 , v52 , v52 , v52 , v52 , v52 , v52 , v52 , v52 , v52 , v52 , v52 , v52 , v52 , v52 , v52 , v52 , v52 , v52 , v52 , v52 , v52 , v52 , v52 , v52 , v52 , v52 , v52 , v52 , v52 , v52 , v52 , v52 , v52 , v52 , v52 , v52 };
wire [63:0] v54 = v53 & v31;
wire [15:0] v55 = 16'b0110111100110100;
wire v56 = v55 == v8;
wire v57 = instruction_bits[17: 17];
wire v58 = v14 == v57;
wire v5a = Advice_3 == v4c;
wire v5b = v5a;
wire v5c = v5b ^ v14;
wire v5d = v14 & v5c & v14;
wire v5e = v56 & v58 & v26 & v5d;
wire v5f = v5e;
wire [63:0] v60 = { v5f , v5f , v5f , v5f , v5f , v5f , v5f , v5f , v5f , v5f , v5f , v5f , v5f , v5f , v5f , v5f , v5f , v5f , v5f , v5f , v5f , v5f , v5f , v5f , v5f , v5f , v5f , v5f , v5f , v5f , v5f , v5f , v5f , v5f , v5f , v5f , v5f , v5f , v5f , v5f , v5f , v5f , v5f , v5f , v5f , v5f , v5f , v5f , v5f , v5f , v5f , v5f , v5f , v5f , v5f , v5f , v5f , v5f , v5f , v5f , v5f , v5f , v5f , v5f };
wire [63:0] v61 = v60 & v1e;
wire [23:0] v62 = 24'b011001000110011010010110;
wire [23:0] v63 = instruction_bits[23: 0];
wire v64 = v62 == v63;
wire [1:0] v65 = 2'b11;
wire [1:0] v66 = instruction_bits[31: 30];
wire v67 = v65 == v66;
wire v68 = v64 & v67 & v41 & v14;
wire v69 = v68;
wire [63:0] v6a = { v69 , v69 , v69 , v69 , v69 , v69 , v69 , v69 , v69 , v69 , v69 , v69 , v69 , v69 , v69 , v69 , v69 , v69 , v69 , v69 , v69 , v69 , v69 , v69 , v69 , v69 , v69 , v69 , v69 , v69 , v69 , v69 , v69 , v69 , v69 , v69 , v69 , v69 , v69 , v69 , v69 , v69 , v69 , v69 , v69 , v69 , v69 , v69 , v69 , v69 , v69 , v69 , v69 , v69 , v69 , v69 , v69 , v69 , v69 , v69 , v69 , v69 , v69 , v69 };
wire [31:0] v6c = 32'b00001000000000000000000000000000;
wire [31:0] v6d = Advice_4 << v6c;
wire [31:0] v6e = v6d >>> v6c;
wire [31:0] pad_111 = (v6e[31:31] == 1'b1) ?32'b11111111111111111111111111111111 : 32'b00000000000000000000000000000000;
wire [63:0] v6f = { pad_111, v6e };
wire [63:0] v70 = v6a & v6f;
wire [23:0] v71 = 24'b011001100110011011101111;
wire v72 = v71 == v63;
wire [4:0] v73 = 5'b10111;
wire [4:0] v74 = instruction_bits[31: 27];
wire v75 = v73 == v74;
wire v76 = v14;
wire v77 = v72 & v75 & vf & v76;
wire v78 = v77;
wire [63:0] v79 = { v78 , v78 , v78 , v78 , v78 , v78 , v78 , v78 , v78 , v78 , v78 , v78 , v78 , v78 , v78 , v78 , v78 , v78 , v78 , v78 , v78 , v78 , v78 , v78 , v78 , v78 , v78 , v78 , v78 , v78 , v78 , v78 , v78 , v78 , v78 , v78 , v78 , v78 , v78 , v78 , v78 , v78 , v78 , v78 , v78 , v78 , v78 , v78 , v78 , v78 , v78 , v78 , v78 , v78 , v78 , v78 , v78 , v78 , v78 , v78 , v78 , v78 , v78 , v78 };
wire [31:0] v7b = Advice_5 << v6c;
wire [31:0] v7c = v7b >>> v6c;
wire [31:0] pad_125 = (v7c[31:31] == 1'b1) ?32'b11111111111111111111111111111111 : 32'b00000000000000000000000000000000;
wire [63:0] v7d = { pad_125, v7c };
wire [63:0] v7e = v79 & v7d;
wire [31:0] v7f = 32'b01100110011001101110111110110100;
wire [31:0] v80 = instruction_bits[31: 0];
wire v81 = v7f == v80;
wire [55:0] v82 = 56'b00000000000000000000000000000000000000000000000000000000;
wire [55:0] v83 = instruction_bits[119: 64];
wire v84 = v82 == v83;
wire v85 = v81 & v84 & v38;
wire v86 = v85;
wire [63:0] v87 = { v86 , v86 , v86 , v86 , v86 , v86 , v86 , v86 , v86 , v86 , v86 , v86 , v86 , v86 , v86 , v86 , v86 , v86 , v86 , v86 , v86 , v86 , v86 , v86 , v86 , v86 , v86 , v86 , v86 , v86 , v86 , v86 , v86 , v86 , v86 , v86 , v86 , v86 , v86 , v86 , v86 , v86 , v86 , v86 , v86 , v86 , v86 , v86 , v86 , v86 , v86 , v86 , v86 , v86 , v86 , v86 , v86 , v86 , v86 , v86 , v86 , v86 , v86 , v86 };
wire [15:0] v88 = v1b[15:0];
wire [15:0] pad_137 = (v88[15:15] == 1'b1) ?16'b1111111111111111 : 16'b0000000000000000;
wire [31:0] v89 = { pad_137, v88 };
wire [31:0] pad_138 = (v89[31:31] == 1'b1) ?32'b11111111111111111111111111111111 : 32'b00000000000000000000000000000000;
wire [63:0] v8a = { pad_138, v89 };
wire [63:0] v8b = v87 & v8a;
wire [15:0] v8c = 16'b0110111100110101;
wire v8d = v8c == v8;
wire v8e = v8d & v37 & v5d;
wire v8f = v8e;
wire [63:0] v90 = { v8f , v8f , v8f , v8f , v8f , v8f , v8f , v8f , v8f , v8f , v8f , v8f , v8f , v8f , v8f , v8f , v8f , v8f , v8f , v8f , v8f , v8f , v8f , v8f , v8f , v8f , v8f , v8f , v8f , v8f , v8f , v8f , v8f , v8f , v8f , v8f , v8f , v8f , v8f , v8f , v8f , v8f , v8f , v8f , v8f , v8f , v8f , v8f , v8f , v8f , v8f , v8f , v8f , v8f , v8f , v8f , v8f , v8f , v8f , v8f , v8f , v8f , v8f , v8f };
wire [63:0] v91 = v90 & v1e;
wire [15:0] v92 = 16'b0110011001101111;
wire v93 = v92 == v8;
wire [4:0] v94 = instruction_bits[23: 19];
wire v95 = v49 == v94;
wire v97 = Advice_6 == v4c;
wire v98 = v97;
wire v99 = v98 ^ v14;
wire v9a = v99 & v14 & v4f;
wire v9b = v93 & v95 & v37 & v9a;
wire v9c = v9b;
wire [63:0] v9d = { v9c , v9c , v9c , v9c , v9c , v9c , v9c , v9c , v9c , v9c , v9c , v9c , v9c , v9c , v9c , v9c , v9c , v9c , v9c , v9c , v9c , v9c , v9c , v9c , v9c , v9c , v9c , v9c , v9c , v9c , v9c , v9c , v9c , v9c , v9c , v9c , v9c , v9c , v9c , v9c , v9c , v9c , v9c , v9c , v9c , v9c , v9c , v9c , v9c , v9c , v9c , v9c , v9c , v9c , v9c , v9c , v9c , v9c , v9c , v9c , v9c , v9c , v9c , v9c };
wire [63:0] v9e = v9d & v31;
wire [15:0] v9f = 16'b0110011010010110;
wire va0 = v9f == v8;
wire [1:0] va1 = instruction_bits[23: 22];
wire va2 = v65 == va1;
wire [79:0] va3 = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
wire [79:0] va4 = instruction_bits[119: 40];
wire va5 = va3 == va4;
wire va6 = va0 & va2 & va5 & v14;
wire va7 = va6;
wire [63:0] va8 = { va7 , va7 , va7 , va7 , va7 , va7 , va7 , va7 , va7 , va7 , va7 , va7 , va7 , va7 , va7 , va7 , va7 , va7 , va7 , va7 , va7 , va7 , va7 , va7 , va7 , va7 , va7 , va7 , va7 , va7 , va7 , va7 , va7 , va7 , va7 , va7 , va7 , va7 , va7 , va7 , va7 , va7 , va7 , va7 , va7 , va7 , va7 , va7 , va7 , va7 , va7 , va7 , va7 , va7 , va7 , va7 , va7 , va7 , va7 , va7 , va7 , va7 , va7 , va7 };
wire [63:0] va9 = va8 & v6f;
wire [23:0] vaa = 24'b101001100010011010010110;
wire vab = vaa == v63;
wire vac = vab & v67 & v84 & v14;
wire [15:0] vad = 16'b0110010011010110;
wire vae = vad == v8;
wire vaf = vae & va2 & vf & v14;
wire [7:0] vb0 = 8'b10010110;
wire vb1 = vb0 == v47;
wire [1:0] vb2 = instruction_bits[15: 14];
wire vb3 = v65 == vb2;
wire vb4 = vb1 & vb3 & v41 & v14;
wire [15:0] vb5 = 16'b1110011010010110;
wire vb6 = vb5 == v8;
wire vb7 = vb6 & va2 & v37 & v14;
wire [23:0] vb8 = 24'b101001101110011011010110;
wire vb9 = vb8 == v63;
wire vba = vb9 & v67 & va5 & v14;
wire [7:0] vbb = 8'b11010110;
wire vbc = vbb == v47;
wire vbd = vbc & vb3 & v26 & v14;
wire vbe = vac | vaf | vb4 | vb7 | vba | vbd;
wire [63:0] vbf = { vbe , vbe , vbe , vbe , vbe , vbe , vbe , vbe , vbe , vbe , vbe , vbe , vbe , vbe , vbe , vbe , vbe , vbe , vbe , vbe , vbe , vbe , vbe , vbe , vbe , vbe , vbe , vbe , vbe , vbe , vbe , vbe , vbe , vbe , vbe , vbe , vbe , vbe , vbe , vbe , vbe , vbe , vbe , vbe , vbe , vbe , vbe , vbe , vbe , vbe , vbe , vbe , vbe , vbe , vbe , vbe , vbe , vbe , vbe , vbe , vbe , vbe , vbe , vbe };
wire [31:0] pad_192 = (Advice_4[31:31] == 1'b1) ?32'b11111111111111111111111111111111 : 32'b00000000000000000000000000000000;
wire [63:0] vc0 = { pad_192, Advice_4 };
wire [63:0] vc1 = vbf & vc0;
wire [15:0] vc2 = 16'b0110110011101111;
wire vc3 = vc2 == v8;
wire [4:0] vc4 = 5'b00111;
wire vc5 = vc4 == v94;
wire vc6 = vc3 & vc5 & v26 & v76;
wire [7:0] vc7 = 8'b11101111;
wire vc8 = vc7 == v47;
wire vc9 = vc4 == v4a;
wire [103:0] vca = 104'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
wire [103:0] vcb = instruction_bits[119: 16];
wire vcc = vca == vcb;
wire vcd = vc8 & vc9 & vcc & v76;
wire vce = vc6 | vcd;
wire [63:0] vcf = { vce , vce , vce , vce , vce , vce , vce , vce , vce , vce , vce , vce , vce , vce , vce , vce , vce , vce , vce , vce , vce , vce , vce , vce , vce , vce , vce , vce , vce , vce , vce , vce , vce , vce , vce , vce , vce , vce , vce , vce , vce , vce , vce , vce , vce , vce , vce , vce , vce , vce , vce , vce , vce , vce , vce , vce , vce , vce , vce , vce , vce , vce , vce , vce };
wire [63:0] vd0 = { 32'b00000000000000000000000000000000, In_register_EAX };
wire [63:0] vd1 = vcf & vd0;
wire [5:0] vd2 = 6'b010100;
wire vd3 = vd2 == vb;
wire vd4 = v9 & vd3 & v26 & v16;
wire vd5 = vd4;
wire [63:0] vd6 = { vd5 , vd5 , vd5 , vd5 , vd5 , vd5 , vd5 , vd5 , vd5 , vd5 , vd5 , vd5 , vd5 , vd5 , vd5 , vd5 , vd5 , vd5 , vd5 , vd5 , vd5 , vd5 , vd5 , vd5 , vd5 , vd5 , vd5 , vd5 , vd5 , vd5 , vd5 , vd5 , vd5 , vd5 , vd5 , vd5 , vd5 , vd5 , vd5 , vd5 , vd5 , vd5 , vd5 , vd5 , vd5 , vd5 , vd5 , vd5 , vd5 , vd5 , vd5 , vd5 , vd5 , vd5 , vd5 , vd5 , vd5 , vd5 , vd5 , vd5 , vd5 , vd5 , vd5 , vd5 };
wire [63:0] vd7 = vd6 & v1e;
wire [1:0] vd8 = 2'b00;
wire vd9 = vd8 == va1;
wire vda = v14 & v14 & v14 & v14;
wire vdb = va0 & v58 & vd9 & va5 & vda;
wire vdc = vdb;
wire [63:0] vdd = { vdc , vdc , vdc , vdc , vdc , vdc , vdc , vdc , vdc , vdc , vdc , vdc , vdc , vdc , vdc , vdc , vdc , vdc , vdc , vdc , vdc , vdc , vdc , vdc , vdc , vdc , vdc , vdc , vdc , vdc , vdc , vdc , vdc , vdc , vdc , vdc , vdc , vdc , vdc , vdc , vdc , vdc , vdc , vdc , vdc , vdc , vdc , vdc , vdc , vdc , vdc , vdc , vdc , vdc , vdc , vdc , vdc , vdc , vdc , vdc , vdc , vdc , vdc , vdc };
wire [63:0] vde = vdd & v6f;
wire [23:0] vdf = 24'b111011110011010010100110;
wire ve0 = vdf == v63;
wire ve1 = ve0 & v37 & v38;
wire [23:0] ve2 = 24'b001001101110111100110101;
wire ve3 = ve2 == v63;
wire ve4 = ve3 & v84 & v5d;
wire ve5 = instruction_bits[9: 9];
wire ve6 = v14 == ve5;
wire [4:0] ve7 = 5'b10110;
wire ve8 = ve7 == v4a;
wire ve9 = vc8 & ve6 & ve8 & v26 & v38;
wire [15:0] vea = 16'b1110111100110110;
wire veb = vea == v8;
wire vec = veb & vc5 & vf & v38;
wire [4:0] ved = 5'b10101;
wire vee = ved == v4a;
wire vef = vc8 & vee & v41 & v9a;
wire [16:0] vf0 = 17'b11100110111011111;
wire [16:0] vf1 = instruction_bits[16: 0];
wire vf2 = vf0 == vf1;
wire [5:0] vf3 = 6'b110100;
wire vf4 = vf3 == vb;
wire vf5 = vf2 & vf4 & v26 & v38;
wire [4:0] vf6 = 5'b10100;
wire vf7 = vf6 == v4a;
wire vf8 = vc8 & vf7 & vcc & v38;
wire [1:0] vf9 = 2'b10;
wire vfa = vf9 == va1;
wire vfc = Advice_7 == v4c;
wire vfd = vfc;
wire vfe = vfd ^ v14;
wire vff = v14 & v5c & v14 & vfe;
wire v100 = vae & vfa & va5 & vff;
wire v101 = vf9 == vb2;
wire v102 = vbc & v101 & vf & vff;
wire [10:0] v103 = 11'b10010110001;
wire [10:0] v104 = instruction_bits[10: 0];
wire v105 = v103 == v104;
wire v106 = vd8 == vb2;
wire v107 = Advice_7 == v28;
wire v108 = v107;
wire v109 = v108 ^ v14;
wire v10a = v14 & v14 & v4f & v109;
wire v10b = v105 & v106 & v37 & v10a;
wire [10:0] v10c = 11'b10010110101;
wire v10d = v10c == v104;
wire [39:0] v10e = 40'b0000000000000000000000000000000000000000;
wire [39:0] v10f = instruction_bits[119: 80];
wire v110 = v10e == v10f;
wire v111 = v10d & v106 & v110 & vda;
wire [15:0] v112 = 16'b1110011011010110;
wire v113 = v112 == v8;
wire v114 = instruction_bits[18: 18];
wire v115 = v11 == v114;
wire [1:0] v116 = 2'b01;
wire v117 = v116 == va1;
wire v119 = Advice_8;
wire v11a = v119 ^ v14;
wire v11b = v14 & v11a & v14 & v14;
wire v11c = v113 & v115 & v117 & v41 & v11b;
wire [10:0] v11d = 11'b11010110001;
wire v11e = v11d == v104;
wire [4:0] v11f = instruction_bits[18: 14];
wire v120 = v49 == v11f;
wire v121 = v11e & v120 & v23 & v84 & vda;
wire v122 = v116 == vb2;
wire v123 = v14 & v14 & v14 & vfe;
wire v124 = vbc & v122 & v37 & v123;
wire [9:0] v125 = 10'b0010100101;
wire [9:0] v126 = instruction_bits[23: 14];
wire v127 = v125 == v126;
wire [31:0] v128 = 32'b00000000000000000000000000000000;
wire [31:0] v129 = instruction_bits[119: 88];
wire v12a = v128 == v129;
wire v12b = v105 & v127 & v12a & vda;
wire [47:0] v12c = 48'b000000000000000000000000000000000000000000000000;
wire [47:0] v12d = instruction_bits[119: 72];
wire v12e = v12c == v12d;
wire v12f = vb6 & v117 & v12e & vda;
wire v130 = vb6 & vfa & v84 & vda;
wire [1:0] v131 = instruction_bits[18: 17];
wire v132 = v116 == v131;
wire v133 = vb6 & v132 & vd9 & v37 & vda;
wire v134 = vb1 & v101 & v37 & vff;
wire v135 = vb1 & ve6 & v122 & v110 & vda;
wire v136 = v14 & v15 & v14 & v14;
wire v137 = vb6 & v115 & vd9 & v37 & v136;
wire [15:0] v138 = 16'b1110111110110100;
wire v139 = v138 == v8;
wire v13a = v139 & v41 & v38;
wire [23:0] v13b = 24'b011011001110111100110110;
wire v13c = v13b == v63;
wire v13d = v13c & va5 & v5d;
wire v13e = v105 & v122 & vc5 & v12a & vda;
wire [10:0] v13f = 11'b11010110101;
wire v140 = v13f == v104;
wire v141 = v140 & v106 & v37 & vda;
wire v142 = v113 & v115 & vd9 & vf & v11b;
wire [15:0] v143 = 16'b1110011011101111;
wire v144 = v143 == v8;
wire [5:0] v145 = 6'b010101;
wire v146 = v145 == vb;
wire v148 = Advice_9;
wire v149 = v148 ^ v14;
wire v14a = v149 & v14 & v14;
wire v14b = v144 & v146 & va5 & v14a;
wire v14c = vae & v58 & vd9 & vf & vda;
wire v14d = v14 & v14 & v4f & v14;
wire v14e = v105 & v101 & v84 & v14d;
wire [18:0] v14f = 19'b0110010011010110001;
wire [18:0] v150 = instruction_bits[18: 0];
wire v151 = v14f == v150;
wire v152 = v151 & v117 & v12e & v14d;
wire v153 = v105 & v101 & vc5 & v84 & vda;
wire [18:0] v154 = 19'b1010011010010110001;
wire v155 = v154 == v150;
wire v156 = Advice_3 == v28;
wire v157 = v156;
wire v158 = v157 ^ v14;
wire v159 = v14 & v158 & v4f & v109;
wire v15a = v155 & vd9 & v84 & v159;
wire v15b = instruction_bits[28: 28];
wire v15c = v14 == v15b;
wire v15d = v155 & vfa & v15c & v12e & vda;
wire v15e = v11e & v106 & vf & v10a;
wire [18:0] v15f = 19'b1010011010010110101;
wire v160 = v15f == v150;
wire v161 = v160 & vd9 & v12a & vda;
wire [2:0] v162 = 3'b000;
wire v163 = Advice_3 == v162;
wire [2:0] v164 = 3'b100;
wire v165 = Advice_3 == v164;
wire [2:0] v166 = 3'b010;
wire v167 = Advice_3 == v166;
wire [2:0] v168 = 3'b110;
wire v169 = Advice_3 == v168;
wire [2:0] v16a = 3'b011;
wire v16b = Advice_3 == v16a;
wire [2:0] v16c = 3'b111;
wire v16d = Advice_3 == v16c;
wire v16e = v163 & v165 & v167 & v169 & v16b & v16d;
wire v16f = v16e ^ v14;
wire v170 = v14 & v16f & v4f & v14;
wire v171 = v11e & v122 & v84 & v170;
wire v172 = vb1 & v106 & v41 & vda;
wire v173 = v105 & v120 & v12a & v14d;
wire v174 = v11e & v101 & va5 & v170;
wire [16:0] v175 = 17'b11100110110101101;
wire v176 = v175 == vf1;
wire v177 = v14 == v114;
wire v178 = v176 & v177 & vd9 & vf & vda;
wire [15:0] v179 = 16'b0010011010010110;
wire v17a = v179 == v8;
wire v17b = v17a & v58 & vfa & v84 & vda;
wire [18:0] v17c = 19'b0010011011010110001;
wire v17d = v17c == v150;
wire v17e = v17d & vfa & v41 & v14d;
wire v17f = v105 & v122 & v12a & v14d;
wire [15:0] v180 = 16'b0110010010010110;
wire v181 = v180 == v8;
wire v182 = v181 & v117 & v12a & vff;
wire v183 = v11e & v122 & vc5 & v84 & vda;
wire v184 = v14 & v14 & v14 & v109;
wire v185 = v11e & v106 & vc5 & vf & v184;
wire v186 = v113 & v115 & vfa & va5 & v11b;
wire v187 = v11e & v101 & vc5 & va5 & vda;
wire [9:0] v188 = 10'b0010100111;
wire v189 = v188 == v126;
wire v18a = v11e & v189 & v84 & vda;
wire [15:0] v18b = 16'b1110111100110100;
wire v18c = v18b == v8;
wire v18d = v18c & v58 & vc5 & v26 & v38;
wire v18e = instruction_bits[25: 25];
wire v18f = v14 == v18e;
wire v190 = v151 & vd9 & v18f & va5 & v14d;
wire [18:0] v191 = 19'b0110110010010110001;
wire v192 = v191 == v150;
wire [23:0] v193 = 24'b000000000000000000000000;
wire [23:0] v194 = instruction_bits[119: 96];
wire v195 = v193 == v194;
wire v196 = v192 & v117 & v195 & v14d;
wire [16:0] v197 = 17'b11100110100101101;
wire v198 = v197 == vf1;
wire v199 = v198 & v177 & vd9 & v37 & vda;
wire v19a = v17a & vd9 & v37 & vda;
wire v19b = Advice_6 == v162;
wire v19c = Advice_6 == v164;
wire v19d = Advice_6 == v166;
wire v19e = Advice_6 == v168;
wire v19f = Advice_6 == v16a;
wire v1a0 = Advice_6 == v16c;
wire v1a1 = v19b & v19c & v19d & v19e & v19f & v1a0;
wire v1a2 = v1a1 ^ v14;
wire v1a3 = v1a2 & v14 & v14;
wire v1a4 = veb & v23 & vf & v1a3;
wire [18:0] v1a5 = 19'b0010011011010110101;
wire v1a6 = v1a5 == v150;
wire v1a7 = v1a6 & vd9 & v84 & vda;
wire v1a8 = vae & v117 & v84 & vff;
wire v1a9 = v105 & v106 & vc5 & v37 & v184;
wire v1aa = vbc & v106 & v26 & vda;
wire v1ab = ve1 | ve4 | ve9 | vec | vef | vf5 | vf8 | v100 | v102 | v10b | v111 | v11c | v121 | v124 | v12b | v12f | v130 | v133 | v134 | v135 | v137 | v13a | v13d | v13e | v141 | v142 | v14b | v14c | v14e | v152 | v153 | v15a | v15d | v15e | v161 | v171 | v172 | v173 | v174 | v178 | v17b | v17e | v17f | v182 | v183 | v185 | v186 | v187 | v18a | v18d | v190 | v196 | v199 | v19a | v1a4 | v1a7 | v1a8 | v1a9 | v1aa;
wire [63:0] v1ac = { v1ab , v1ab , v1ab , v1ab , v1ab , v1ab , v1ab , v1ab , v1ab , v1ab , v1ab , v1ab , v1ab , v1ab , v1ab , v1ab , v1ab , v1ab , v1ab , v1ab , v1ab , v1ab , v1ab , v1ab , v1ab , v1ab , v1ab , v1ab , v1ab , v1ab , v1ab , v1ab , v1ab , v1ab , v1ab , v1ab , v1ab , v1ab , v1ab , v1ab , v1ab , v1ab , v1ab , v1ab , v1ab , v1ab , v1ab , v1ab , v1ab , v1ab , v1ab , v1ab , v1ab , v1ab , v1ab , v1ab , v1ab , v1ab , v1ab , v1ab , v1ab , v1ab , v1ab , v1ab };
wire [31:0] pad_429 = (v1b[31:31] == 1'b1) ?32'b11111111111111111111111111111111 : 32'b00000000000000000000000000000000;
wire [63:0] v1ad = { pad_429, v1b };
wire [63:0] v1ae = v1ac & v1ad;
wire [18:0] v1af = 19'b0110011010010110001;
wire v1b0 = v1af == v150;
wire v1b1 = v1b0 & vfa & v37 & v14d;
wire v1b2 = v1b1;
wire [63:0] v1b3 = { v1b2 , v1b2 , v1b2 , v1b2 , v1b2 , v1b2 , v1b2 , v1b2 , v1b2 , v1b2 , v1b2 , v1b2 , v1b2 , v1b2 , v1b2 , v1b2 , v1b2 , v1b2 , v1b2 , v1b2 , v1b2 , v1b2 , v1b2 , v1b2 , v1b2 , v1b2 , v1b2 , v1b2 , v1b2 , v1b2 , v1b2 , v1b2 , v1b2 , v1b2 , v1b2 , v1b2 , v1b2 , v1b2 , v1b2 , v1b2 , v1b2 , v1b2 , v1b2 , v1b2 , v1b2 , v1b2 , v1b2 , v1b2 , v1b2 , v1b2 , v1b2 , v1b2 , v1b2 , v1b2 , v1b2 , v1b2 , v1b2 , v1b2 , v1b2 , v1b2 , v1b2 , v1b2 , v1b2 , v1b2 };
wire [63:0] v1b4 = v1b3 & v6f;
wire v1b5 = v1b0 & v117 & v110 & v14d;
wire v1b6 = v1b5;
wire [63:0] v1b7 = { v1b6 , v1b6 , v1b6 , v1b6 , v1b6 , v1b6 , v1b6 , v1b6 , v1b6 , v1b6 , v1b6 , v1b6 , v1b6 , v1b6 , v1b6 , v1b6 , v1b6 , v1b6 , v1b6 , v1b6 , v1b6 , v1b6 , v1b6 , v1b6 , v1b6 , v1b6 , v1b6 , v1b6 , v1b6 , v1b6 , v1b6 , v1b6 , v1b6 , v1b6 , v1b6 , v1b6 , v1b6 , v1b6 , v1b6 , v1b6 , v1b6 , v1b6 , v1b6 , v1b6 , v1b6 , v1b6 , v1b6 , v1b6 , v1b6 , v1b6 , v1b6 , v1b6 , v1b6 , v1b6 , v1b6 , v1b6 , v1b6 , v1b6 , v1b6 , v1b6 , v1b6 , v1b6 , v1b6 , v1b6 };
wire [63:0] v1b8 = v1b7 & v6f;
wire [15:0] v1b9 = 16'b1110111100100110;
wire v1ba = v1b9 == v8;
wire v1bb = v1ba & vf & v5d;
wire v1bc = v1ba & v95 & vf & v38;
wire [23:0] v1bd = 24'b011001001110111100100101;
wire v1be = v1bd == v63;
wire v1bf = v1be & v84 & v5d;
wire [23:0] v1c0 = 24'b101001101110111100100110;
wire v1c1 = v1c0 == v63;
wire v1c2 = v1c1 & va5 & v5d;
wire [15:0] v1c3 = 16'b1110111100100100;
wire v1c4 = v1c3 == v8;
wire v1c5 = Advice_6 == v28;
wire v1c6 = v1c5;
wire v1c7 = v1c6 ^ v14;
wire v1c8 = v1c7 & v14 & v2b;
wire v1c9 = v1c4 & vc5 & v26 & v1c8;
wire [4:0] v1ca = 5'b00100;
wire v1cb = v1ca == v4a;
wire v1cc = vc8 & v1cb & vcc & v38;
wire [4:0] v1cd = 5'b00110;
wire v1ce = v1cd == v4a;
wire v1cf = vc8 & ve6 & v1ce & v26 & v38;
wire v1d0 = v1bb | v1bc | v1bf | v1c2 | v1c9 | v1cc | v1cf;
wire [63:0] v1d1 = { v1d0 , v1d0 , v1d0 , v1d0 , v1d0 , v1d0 , v1d0 , v1d0 , v1d0 , v1d0 , v1d0 , v1d0 , v1d0 , v1d0 , v1d0 , v1d0 , v1d0 , v1d0 , v1d0 , v1d0 , v1d0 , v1d0 , v1d0 , v1d0 , v1d0 , v1d0 , v1d0 , v1d0 , v1d0 , v1d0 , v1d0 , v1d0 , v1d0 , v1d0 , v1d0 , v1d0 , v1d0 , v1d0 , v1d0 , v1d0 , v1d0 , v1d0 , v1d0 , v1d0 , v1d0 , v1d0 , v1d0 , v1d0 , v1d0 , v1d0 , v1d0 , v1d0 , v1d0 , v1d0 , v1d0 , v1d0 , v1d0 , v1d0 , v1d0 , v1d0 , v1d0 , v1d0 , v1d0 , v1d0 };
wire [63:0] v1d2 = { 32'b00000000000000000000000000000000, v1b };
wire [63:0] v1d3 = v1d1 & v1d2;
wire [23:0] v1d4 = 24'b011001100110111100100100;
wire v1d5 = v1d4 == v63;
wire v1d6 = v1d5 & v18f & vf & v5d;
wire v1d7 = v1d6;
wire [63:0] v1d8 = { v1d7 , v1d7 , v1d7 , v1d7 , v1d7 , v1d7 , v1d7 , v1d7 , v1d7 , v1d7 , v1d7 , v1d7 , v1d7 , v1d7 , v1d7 , v1d7 , v1d7 , v1d7 , v1d7 , v1d7 , v1d7 , v1d7 , v1d7 , v1d7 , v1d7 , v1d7 , v1d7 , v1d7 , v1d7 , v1d7 , v1d7 , v1d7 , v1d7 , v1d7 , v1d7 , v1d7 , v1d7 , v1d7 , v1d7 , v1d7 , v1d7 , v1d7 , v1d7 , v1d7 , v1d7 , v1d7 , v1d7 , v1d7 , v1d7 , v1d7 , v1d7 , v1d7 , v1d7 , v1d7 , v1d7 , v1d7 , v1d7 , v1d7 , v1d7 , v1d7 , v1d7 , v1d7 , v1d7 , v1d7 };
wire [63:0] v1d9 = v1d8 & v31;
wire v1da = v1cd == v74;
wire v1db = v14 & v158 & v14 & v109;
wire v1dc = v1b0 & vd9 & v1da & v41 & v1db;
wire v1dd = v1dc;
wire [63:0] v1de = { v1dd , v1dd , v1dd , v1dd , v1dd , v1dd , v1dd , v1dd , v1dd , v1dd , v1dd , v1dd , v1dd , v1dd , v1dd , v1dd , v1dd , v1dd , v1dd , v1dd , v1dd , v1dd , v1dd , v1dd , v1dd , v1dd , v1dd , v1dd , v1dd , v1dd , v1dd , v1dd , v1dd , v1dd , v1dd , v1dd , v1dd , v1dd , v1dd , v1dd , v1dd , v1dd , v1dd , v1dd , v1dd , v1dd , v1dd , v1dd , v1dd , v1dd , v1dd , v1dd , v1dd , v1dd , v1dd , v1dd , v1dd , v1dd , v1dd , v1dd , v1dd , v1dd , v1dd , v1dd };
wire [63:0] v1df = v1de & v6f;
wire [15:0] v1e0 = 16'b0110010001101111;
wire v1e1 = v1e0 == v8;
wire v1e2 = ved == v94;
wire v1e3 = v1e1 & v1e2 & v37 & v9a;
wire v1e4 = v1e3;
wire [63:0] v1e5 = { v1e4 , v1e4 , v1e4 , v1e4 , v1e4 , v1e4 , v1e4 , v1e4 , v1e4 , v1e4 , v1e4 , v1e4 , v1e4 , v1e4 , v1e4 , v1e4 , v1e4 , v1e4 , v1e4 , v1e4 , v1e4 , v1e4 , v1e4 , v1e4 , v1e4 , v1e4 , v1e4 , v1e4 , v1e4 , v1e4 , v1e4 , v1e4 , v1e4 , v1e4 , v1e4 , v1e4 , v1e4 , v1e4 , v1e4 , v1e4 , v1e4 , v1e4 , v1e4 , v1e4 , v1e4 , v1e4 , v1e4 , v1e4 , v1e4 , v1e4 , v1e4 , v1e4 , v1e4 , v1e4 , v1e4 , v1e4 , v1e4 , v1e4 , v1e4 , v1e4 , v1e4 , v1e4 , v1e4 , v1e4 };
wire [63:0] v1e6 = v1e5 & v1e;
wire [18:0] v1e7 = 19'b0110111100100100101;
wire v1e8 = v1e7 == v150;
wire v1e9 = v1e8 & v37 & v5d;
wire v1ea = v1e9;
wire [63:0] v1eb = { v1ea , v1ea , v1ea , v1ea , v1ea , v1ea , v1ea , v1ea , v1ea , v1ea , v1ea , v1ea , v1ea , v1ea , v1ea , v1ea , v1ea , v1ea , v1ea , v1ea , v1ea , v1ea , v1ea , v1ea , v1ea , v1ea , v1ea , v1ea , v1ea , v1ea , v1ea , v1ea , v1ea , v1ea , v1ea , v1ea , v1ea , v1ea , v1ea , v1ea , v1ea , v1ea , v1ea , v1ea , v1ea , v1ea , v1ea , v1ea , v1ea , v1ea , v1ea , v1ea , v1ea , v1ea , v1ea , v1ea , v1ea , v1ea , v1ea , v1ea , v1ea , v1ea , v1ea , v1ea };
wire [63:0] v1ec = v1eb & v31;
wire [18:0] v1ed = 19'b0110111100110100101;
wire v1ee = v1ed == v150;
wire v1ef = v1ee & v37 & v5d;
wire v1f0 = v1ef;
wire [63:0] v1f1 = { v1f0 , v1f0 , v1f0 , v1f0 , v1f0 , v1f0 , v1f0 , v1f0 , v1f0 , v1f0 , v1f0 , v1f0 , v1f0 , v1f0 , v1f0 , v1f0 , v1f0 , v1f0 , v1f0 , v1f0 , v1f0 , v1f0 , v1f0 , v1f0 , v1f0 , v1f0 , v1f0 , v1f0 , v1f0 , v1f0 , v1f0 , v1f0 , v1f0 , v1f0 , v1f0 , v1f0 , v1f0 , v1f0 , v1f0 , v1f0 , v1f0 , v1f0 , v1f0 , v1f0 , v1f0 , v1f0 , v1f0 , v1f0 , v1f0 , v1f0 , v1f0 , v1f0 , v1f0 , v1f0 , v1f0 , v1f0 , v1f0 , v1f0 , v1f0 , v1f0 , v1f0 , v1f0 , v1f0 , v1f0 };
wire [63:0] v1f2 = v1f1 & v1e;
wire v1f3 = va0 & v117 & v12e & vff;
wire v1f4 = v1f3;
wire [63:0] v1f5 = { v1f4 , v1f4 , v1f4 , v1f4 , v1f4 , v1f4 , v1f4 , v1f4 , v1f4 , v1f4 , v1f4 , v1f4 , v1f4 , v1f4 , v1f4 , v1f4 , v1f4 , v1f4 , v1f4 , v1f4 , v1f4 , v1f4 , v1f4 , v1f4 , v1f4 , v1f4 , v1f4 , v1f4 , v1f4 , v1f4 , v1f4 , v1f4 , v1f4 , v1f4 , v1f4 , v1f4 , v1f4 , v1f4 , v1f4 , v1f4 , v1f4 , v1f4 , v1f4 , v1f4 , v1f4 , v1f4 , v1f4 , v1f4 , v1f4 , v1f4 , v1f4 , v1f4 , v1f4 , v1f4 , v1f4 , v1f4 , v1f4 , v1f4 , v1f4 , v1f4 , v1f4 , v1f4 , v1f4 , v1f4 };
wire [63:0] v1f6 = v1f5 & v6f;
wire v1f7 = v73 == v4a;
wire v1f8 = vc8 & v1f7 & vcc & v76;
wire v1f9 = v73 == v94;
wire v1fa = v144 & v1f9 & v26 & v76;
wire v1fb = v1f8 | v1fa;
wire [63:0] v1fc = { v1fb , v1fb , v1fb , v1fb , v1fb , v1fb , v1fb , v1fb , v1fb , v1fb , v1fb , v1fb , v1fb , v1fb , v1fb , v1fb , v1fb , v1fb , v1fb , v1fb , v1fb , v1fb , v1fb , v1fb , v1fb , v1fb , v1fb , v1fb , v1fb , v1fb , v1fb , v1fb , v1fb , v1fb , v1fb , v1fb , v1fb , v1fb , v1fb , v1fb , v1fb , v1fb , v1fb , v1fb , v1fb , v1fb , v1fb , v1fb , v1fb , v1fb , v1fb , v1fb , v1fb , v1fb , v1fb , v1fb , v1fb , v1fb , v1fb , v1fb , v1fb , v1fb , v1fb , v1fb };
wire [31:0] pad_509 = (In_register_EAX[31:31] == 1'b1) ?32'b11111111111111111111111111111111 : 32'b00000000000000000000000000000000;
wire [63:0] v1fd = { pad_509, In_register_EAX };
wire [63:0] v1fe = v1fc & v1fd;
wire [23:0] v1ff = 24'b011001101110111100110100;
wire v200 = v1ff == v63;
wire v201 = v200 & v18f & vf & v5d;
wire v202 = v201;
wire [63:0] v203 = { v202 , v202 , v202 , v202 , v202 , v202 , v202 , v202 , v202 , v202 , v202 , v202 , v202 , v202 , v202 , v202 , v202 , v202 , v202 , v202 , v202 , v202 , v202 , v202 , v202 , v202 , v202 , v202 , v202 , v202 , v202 , v202 , v202 , v202 , v202 , v202 , v202 , v202 , v202 , v202 , v202 , v202 , v202 , v202 , v202 , v202 , v202 , v202 , v202 , v202 , v202 , v202 , v202 , v202 , v202 , v202 , v202 , v202 , v202 , v202 , v202 , v202 , v202 , v202 };
wire [63:0] v204 = v203 & v8a;
wire v205 = va0 & vfa & v41 & v123;
wire v206 = v205;
wire [63:0] v207 = { v206 , v206 , v206 , v206 , v206 , v206 , v206 , v206 , v206 , v206 , v206 , v206 , v206 , v206 , v206 , v206 , v206 , v206 , v206 , v206 , v206 , v206 , v206 , v206 , v206 , v206 , v206 , v206 , v206 , v206 , v206 , v206 , v206 , v206 , v206 , v206 , v206 , v206 , v206 , v206 , v206 , v206 , v206 , v206 , v206 , v206 , v206 , v206 , v206 , v206 , v206 , v206 , v206 , v206 , v206 , v206 , v206 , v206 , v206 , v206 , v206 , v206 , v206 , v206 };
wire [63:0] v208 = v207 & v6f;
wire v209 = v1f | v32 | v3c | v45 | v54 | v61 | v70 | v7e | v8b | v91 | v9e | va9 | vc1 | vd1 | vd7 | vde | v1ae | v1b4 | v1b8 | v1d3 | v1d9 | v1df | v1e6 | v1ec | v1f2 | v1f6 | v1fe | v204 | v208;
wire [7:0] v20a = In_register_EAX[7:0];
wire [7:0] pad_523 = (v20a[7:7] == 1'b1) ?8'b11111111 : 8'b00000000;
wire [15:0] v20b = { pad_523, v20a };
wire [15:0] pad_524 = (v20b[15:15] == 1'b1) ?48'b111111111111111111111111111111111111111111111111 : 48'b000000000000000000000000000000000000000000000000;
wire [63:0] v20c = { pad_524, v20b };
wire [63:0] v20d = v1f1 & v20c;
wire [63:0] v20e = v19 & v20c;
wire [63:0] v20f = v90 & v20c;
wire [63:0] v210 = v1e5 & v20c;
wire [63:0] v211 = vd6 & v20c;
wire [15:0] v212 = { 8'b00000000, v20a };
wire [15:0] pad_531 = (v212[15:15] == 1'b1) ?48'b111111111111111111111111111111111111111111111111 : 48'b000000000000000000000000000000000000000000000000;
wire [63:0] v213 = { pad_531, v212 };
wire [63:0] v214 = v1d8 & v213;
wire v215 = ve4 | ve9 | ve1 | vf8 | v13d | v14b | v18d | v13a | vec | v1a4 | vef | vf5;
wire [63:0] v216 = { v215 , v215 , v215 , v215 , v215 , v215 , v215 , v215 , v215 , v215 , v215 , v215 , v215 , v215 , v215 , v215 , v215 , v215 , v215 , v215 , v215 , v215 , v215 , v215 , v215 , v215 , v215 , v215 , v215 , v215 , v215 , v215 , v215 , v215 , v215 , v215 , v215 , v215 , v215 , v215 , v215 , v215 , v215 , v215 , v215 , v215 , v215 , v215 , v215 , v215 , v215 , v215 , v215 , v215 , v215 , v215 , v215 , v215 , v215 , v215 , v215 , v215 , v215 , v215 };
wire [63:0] v217 = v216 & v1fd;
wire [63:0] v218 = v44 & v213;
wire [63:0] v219 = v2f & v213;
wire [63:0] v21a = v53 & v213;
wire [15:0] v21b = In_register_EAX[15:0];
wire [15:0] pad_540 = (v21b[15:15] == 1'b1) ?16'b1111111111111111 : 16'b0000000000000000;
wire [31:0] v21c = { pad_540, v21b };
wire [31:0] pad_541 = (v21c[31:31] == 1'b1) ?32'b11111111111111111111111111111111 : 32'b00000000000000000000000000000000;
wire [63:0] v21d = { pad_541, v21c };
wire [63:0] v21e = v203 & v21d;
wire [63:0] v21f = vdd & v8a;
wire [63:0] v220 = v207 & v8a;
wire [63:0] v221 = v9d & v213;
wire [63:0] v222 = v87 & v21d;
wire [63:0] v223 = v60 & v20c;
wire v224 = v100 | v10b | v111 | v11c | v124 | v12f | v130 | v133 | v134 | v135 | v137 | v13e | v142 | v12b | v14e | v102 | v152 | v153 | v15a | v15e | v171 | v172 | v161 | v173 | v174 | v178 | v17e | v182 | v183 | v186 | v187 | v18a | v190 | v196 | v185 | v199 | v19a | v141 | v17b | v17f | v121 | v1a7 | v15d | v1a8 | v14c | v1a9 | v1aa;
wire [63:0] v225 = { v224 , v224 , v224 , v224 , v224 , v224 , v224 , v224 , v224 , v224 , v224 , v224 , v224 , v224 , v224 , v224 , v224 , v224 , v224 , v224 , v224 , v224 , v224 , v224 , v224 , v224 , v224 , v224 , v224 , v224 , v224 , v224 , v224 , v224 , v224 , v224 , v224 , v224 , v224 , v224 , v224 , v224 , v224 , v224 , v224 , v224 , v224 , v224 , v224 , v224 , v224 , v224 , v224 , v224 , v224 , v224 , v224 , v224 , v224 , v224 , v224 , v224 , v224 , v224 };
wire [63:0] v226 = v225 & vc0;
wire [63:0] v227 = { 32'b00000000000000000000000000000000, Advice_5 };
wire [63:0] v228 = vcf & v227;
wire [63:0] v229 = v3b & v213;
wire [63:0] v22a = v1b3 & v8a;
wire [31:0] pad_556 = (Advice_10[31:31] == 1'b1) ?32'b11111111111111111111111111111111 : 32'b00000000000000000000000000000000;
wire [63:0] v22c = { pad_556, Advice_10 };
wire [63:0] v22d = vbf & v22c;
wire [63:0] v22e = v79 & v21d;
wire [31:0] pad_559 = (Advice_5[31:31] == 1'b1) ?32'b11111111111111111111111111111111 : 32'b00000000000000000000000000000000;
wire [63:0] v22f = { pad_559, Advice_5 };
wire [63:0] v230 = v1fc & v22f;
wire [31:0] v231 = Advice_10 << v6c;
wire [31:0] v232 = v231 >>> v6c;
wire [31:0] pad_563 = (v232[31:31] == 1'b1) ?32'b11111111111111111111111111111111 : 32'b00000000000000000000000000000000;
wire [63:0] v233 = { pad_563, v232 };
wire [63:0] v234 = va8 & v233;
wire [63:0] v235 = v6a & v233;
wire [63:0] v236 = v1b7 & v8a;
wire [63:0] v237 = v1eb & v213;
wire [63:0] v238 = v1d1 & vd0;
wire [63:0] v239 = v1f5 & v8a;
wire [63:0] v23a = v1de & v8a;
wire v23b = v20d | v20e | v20f | v210 | v211 | v214 | v217 | v218 | v219 | v21a | v21e | v21f | v220 | v221 | v222 | v223 | v226 | v228 | v229 | v22a | v22d | v22e | v230 | v234 | v235 | v236 | v237 | v238 | v239 | v23a;
wire [63:0] v23c = v209 * v23b;
wire [31:0] v23d = v23c[31:0];
wire [15:0] v23e = v23d[15:0];
wire [31:0] v23f = { 16'b0000000000000000, v23e };
wire [31:0] v240 = v5 | v23f;
wire v242 = v240 == Out_register_EAX;
wire v245 = In_register_EBX == Out_register_EBX;
wire v248 = In_register_ECX == Out_register_ECX;
wire [31:0] v24a = In_register_EDX & v4;
wire [31:0] v24b = v23d >> v6c;
wire [15:0] v24c = v24b[15:0];
wire [31:0] v24d = { 16'b0000000000000000, v24c };
wire [31:0] v24e = v24a | v24d;
wire v250 = v24e == Out_register_EDX;
wire v253 = In_register_ESI == Out_register_ESI;
wire v256 = In_register_EDI == Out_register_EDI;
wire v259 = In_register_ESP == Out_register_ESP;
wire v25c = In_register_EBP == Out_register_EBP;
wire [31:0] v25e = 32'b00010000000000000000000000000000;
wire [31:0] v25f = In_register_EIP + v25e;
wire v261 = v25f == Out_register_EIP;
wire v264 = In_register_CSBASE == Out_register_CSBASE;
wire v267 = In_register_SSBASE == Out_register_SSBASE;
wire v26a = In_register_ESBASE == Out_register_ESBASE;
wire v26d = In_register_DSBASE == Out_register_DSBASE;
wire v270 = In_register_GSBASE == Out_register_GSBASE;
wire v273 = In_register_FSBASE == Out_register_FSBASE;
wire v276 = In_register_AF == Out_register_AF;
wire [31:0] v277 = 32'b00000000000000011111111111111111;
wire [31:0] v278 = v23d + v277;
wire v279 = v278 < v4;
wire v27b = v279 == Out_register_CF;
wire v27e = In_register_DF == Out_register_DF;
wire v280 = v279 == Out_register_OF;
wire v283 = In_register_PF == Out_register_PF;
wire v286 = In_register_SF == Out_register_SF;
wire v289 = In_register_ZF == Out_register_ZF;
wire v28a = v242 & v245 & v248 & v250 & v253 & v256 & v259 & v25c & v261 & v264 & v267 & v26a & v26d & v270 & v273 & v276 & v27b & v27e & v280 & v283 & v286 & v289;
wire [31:0] v28c = In_register_DSBASE + v128;
wire [31:0] v28d = v128 << v128;
wire [31:0] v28e = v28c + v28d;
wire [31:0] v28f = instruction_bits[63: 32];
wire [31:0] v291 = v28e + v28f;
wire v292 = v291 == Advice_5;
wire v294 = v11 == Out_error_flag;
wire [3:0] v295 = 4'b0100;
wire v297 =  v295 == memory_0[15: 12] && Advice_5 == memory_0[79: 16] && In_timestamp == memory_0[207: 144] && 4'd0 == memory_0[11: 8] && 1'b1 == memory_0[0: 0] && 6'b000000 == memory_0[7: 2] && 1'b0 == memory_0[1: 1];
wire v299 = In_error_flag == v11;
wire [63:0] v29a = 64'b1000000000000000000000000000000000000000000000000000000000000000;
wire [63:0] v29b = In_timestamp + v29a;
wire v29d = v29b == Out_timestamp;
wire v29e = In_error_flag ^ v14;
wire v29f = v29e | Out_error_flag;
wire v2a0 = v28a & v292 & v294 & v297 & v299 & v85 & v29d & v29f;
wire rnx2x0 = 1'b0 || v2a0;
wire onx2x0 = 1'b0 || ( 1'b0 && v2a0);
wire [31:0] v2a1 = instruction_bits[47: 16];
wire [31:0] v2a3 = v28e + v2a1;
wire v2a4 = v2a3 == Advice_5;
wire v2a5 = v23d == Out_register_EAX;
wire [63:0] v2a6 = 64'b0000010000000000000000000000000000000000000000000000000000000000;
wire [63:0] v2a7 = v23c >> v2a6;
wire [31:0] v2a8 = v2a7[31:0];
wire v2a9 = v2a8 == Out_register_EDX;
wire [31:0] v2aa = 32'b01100000000000000000000000000000;
wire [31:0] v2ab = In_register_EIP + v2aa;
wire v2ac = v2ab == Out_register_EIP;
wire [63:0] v2ad = 64'b0000000000000000000000000000000111111111111111111111111111111111;
wire [63:0] v2ae = v23c + v2ad;
wire [63:0] v2af = 64'b0000000000000000000000000000000011111111111111111111111111111111;
wire v2b0 = v2ae < v2af;
wire v2b1 = v2b0 == Out_register_CF;
wire v2b2 = v2b0 == Out_register_OF;
wire v2b3 = v2a5 & v245 & v248 & v2a9 & v253 & v256 & v259 & v25c & v2ac & v264 & v267 & v26a & v26d & v270 & v273 & v276 & v2b1 & v27e & v2b2 & v283 & v286 & v289;
wire [3:0] v2b4 = 4'b0010;
wire v2b5 =  v2b4 == memory_0[15: 12] && Advice_5 == memory_0[79: 16] && In_timestamp == memory_0[207: 144] && 4'd0 == memory_0[11: 8] && 1'b1 == memory_0[0: 0] && 6'b000000 == memory_0[7: 2] && 1'b0 == memory_0[1: 1];
wire v2b6 = v2a4 & v2b3 & v294 & v13a & v299 & v29f & v2b5 & v29d;
wire rnx2x1 = rnx2x0 || v2b6;
wire onx2x1 = onx2x0 || ( rnx2x0 && v2b6);
wire [31:0] v2b7 = 32'b11100000000000000000000000000000;
wire [31:0] v2b8 = In_register_EIP + v2b7;
wire v2b9 = v2b8 == Out_register_EIP;
wire v2ba = v2a5 & v245 & v248 & v2a9 & v253 & v256 & v259 & v25c & v2b9 & v264 & v267 & v26a & v26d & v270 & v273 & v276 & v2b1 & v27e & v2b2 & v283 & v286 & v289;
wire [31:0] v2bb = instruction_bits[55: 24];
wire [31:0] v2bd = v28e + v2bb;
wire v2be = v2bd == Advice_5;
wire v2bf = v2ba & v2be & v294 & v29d & v299 & v2b5 & ve1 & v29f;
wire rnx2x2 = rnx2x1 || v2bf;
wire onx2x2 = onx2x1 || ( rnx2x1 && v2bf);
wire [31:0] v2c0 = 32'b00000000111111111111111111111111;
wire [31:0] v2c1 = In_register_EAX & v2c0;
wire [15:0] v2c2 = v23c[15:0];
wire [7:0] v2c3 = v2c2[7:0];
wire [31:0] v2c4 = { 24'b000000000000000000000000, v2c3 };
wire [31:0] v2c5 = v2c1 | v2c4;
wire [31:0] v2c6 = 32'b11111111000000001111111111111111;
wire [31:0] v2c7 = v2c5 & v2c6;
wire [15:0] v2c8 = 16'b0001000000000000;
wire [15:0] v2c9 = v2c2 >> v2c8;
wire [7:0] v2ca = v2c9[7:0];
wire [31:0] v2cb = { 24'b000000000000000000000000, v2ca };
wire [31:0] v2cc = v2cb << v25e;
wire [31:0] v2cd = v2c7 | v2cc;
wire v2ce = v2cd == Out_register_EAX;
wire v2cf = In_register_EDX == Out_register_EDX;
wire [15:0] v2d0 = 16'b1111111100000000;
wire v2d1 = v2c2 > v2d0;
wire v2d2 = v2d1 == Out_register_CF;
wire v2d3 = v2d1 == Out_register_OF;
wire v2d4 = v2ce & v245 & v248 & v2cf & v253 & v256 & v259 & v25c & v2ac & v264 & v267 & v26a & v26d & v270 & v273 & v276 & v2d2 & v27e & v2d3 & v283 & v286 & v289;
wire [3:0] v2d5 = 4'b1000;
wire v2d6 =  v2d5 == memory_0[15: 12] && Advice_5 == memory_0[79: 16] && In_timestamp == memory_0[207: 144] && 4'd0 == memory_0[11: 8] && 1'b1 == memory_0[0: 0] && 6'b000000 == memory_0[7: 2] && 1'b0 == memory_0[1: 1];
wire v2d7 = v2a4 & v294 & v2d4 & v29d & v2d6 & v42 & v299 & v29f;
wire rnx2x3 = rnx2x2 || v2d7;
wire onx2x3 = onx2x2 || ( rnx2x2 && v2d7);
wire [31:0] v2d8 = 32'b00100000000000000000000000000000;
wire [31:0] v2d9 = In_register_EIP + v2d8;
wire v2da = v2d9 == Out_register_EIP;
wire v2db = v242 & v245 & v248 & v250 & v253 & v256 & v259 & v25c & v2da & v264 & v267 & v26a & v26d & v270 & v273 & v276 & v27b & v27e & v280 & v283 & v286 & v289;
wire [31:0] v2dd = ( Advice_11 == 3'd0) ? In_register_EAX :
	( Advice_11 == 3'd1) ? In_register_ECX :
	( Advice_11 == 3'd2) ? In_register_EDX :
	( Advice_11 == 3'd3) ? In_register_EBX :
	( Advice_11 == 3'd4) ? In_register_ESP :
	( Advice_11 == 3'd5) ? In_register_EBP :
	( Advice_11 == 3'd6) ? In_register_ESI : In_register_EDI;
wire [31:0] v2de = 32'b11111111111111110000000000000000;
wire [31:0] v2df = v2dd & v2de;
wire v2e0 = v2df == Advice_5;
wire [2:0] v2e1 = instruction_bits[26: 24];
wire [2:0] v2e2 = { v2e1 };
wire v2e3 = v2e2 == Advice_6;
wire v2e4 = Advice_6 == Advice_11;
wire v2e5 = v2db & v2e0 & v294 & v2e3 & v299 & v29f & v77 & v29d & v2e4;
wire rnx2x4 = rnx2x3 || v2e5;
wire onx2x4 = onx2x3 || ( rnx2x3 && v2e5);
wire [31:0] v2e6 = 32'b01000000000000000000000000000000;
wire [31:0] v2e7 = In_register_EIP + v2e6;
wire v2e8 = v2e7 == Out_register_EIP;
wire v2e9 = v2a5 & v245 & v248 & v2a9 & v253 & v256 & v259 & v25c & v2e8 & v264 & v267 & v26a & v26d & v270 & v273 & v276 & v2b1 & v27e & v2b2 & v283 & v286 & v289;
wire v2ea = v2dd == Advice_5;
wire [2:0] v2eb = instruction_bits[10: 8];
wire [2:0] v2ec = { v2eb };
wire v2ed = v2ec == Advice_6;
wire v2ee = v2e9 & v2ea & v294 & v299 & v2ed & v29f & v1f8 & v29d & v2e4;
wire rnx2x5 = rnx2x4 || v2ee;
wire onx2x5 = onx2x4 || ( rnx2x4 && v2ee);
wire [2:0] v2ef = instruction_bits[18: 16];
wire [2:0] v2f0 = { v2ef };
wire v2f1 = v2f0 == Advice_6;
wire [31:0] v2f2 = 32'b11000000000000000000000000000000;
wire [31:0] v2f3 = In_register_EIP + v2f2;
wire v2f4 = v2f3 == Out_register_EIP;
wire v2f5 = v2a5 & v245 & v248 & v2a9 & v253 & v256 & v259 & v25c & v2f4 & v264 & v267 & v26a & v26d & v270 & v273 & v276 & v2b1 & v27e & v2b2 & v283 & v286 & v289;
wire v2f6 = v294 & v299 & v2f1 & v2f5 & v1fa & v2ea & v29d & v29f & v2e4;
wire rnx2x6 = rnx2x5 || v2f6;
wire onx2x6 = onx2x5 || ( rnx2x5 && v2f6);
wire [31:0] v2f7 = { v23d };
wire [31:0] v2f9 = ( Advice_12 == 3'd0) ? Out_register_EAX :
	( Advice_12 == 3'd1) ? Out_register_ECX :
	( Advice_12 == 3'd2) ? Out_register_EDX :
	( Advice_12 == 3'd3) ? Out_register_EBX :
	( Advice_12 == 3'd4) ? Out_register_ESP :
	( Advice_12 == 3'd5) ? Out_register_EBP :
	( Advice_12 == 3'd6) ? Out_register_ESI : Out_register_EDI;
wire v2fa = v2f7 == v2f9;
wire v2fb = In_register_EAX == Out_register_EAX;
wire v2fc = v19b | v2fb;
wire v2fd = v19e | v245;
wire v2fe = v19c | v248;
wire v2ff = v19d | v2cf;
wire v300 = v19f | v253;
wire v301 = v1a0 | v256;
wire v302 = v97 | v259;
wire v303 = v1c5 | v25c;
wire v304 = v2fc & v2fd & v2fe & v2ff & v300 & v301 & v302 & v303 & v2f4 & v264 & v267 & v26a & v26d & v270 & v273 & v276 & v2b1 & v27e & v2b2 & v283 & v286 & v289;
wire v305 = v2fa & v304;
wire v306 = v2dd == Advice_10;
wire v307 = v2ec == Advice_3;
wire [2:0] v308 = instruction_bits[13: 11];
wire [2:0] v309 = { v308 };
wire v30a = v309 == Advice_6;
wire [7:0] v30b = instruction_bits[23: 16];
wire [7:0] pad_780 = (v30b[7:7] == 1'b1) ?24'b111111111111111111111111 : 24'b000000000000000000000000;
wire [31:0] v30c = { pad_780, v30b };
wire v30e = v30c == Advice_4;
wire v30f = Advice_3 == Advice_11;
wire v310 = Advice_6 == Advice_12;
wire v311 = v305 & v306 & v294 & v299 & v307 & v29d & v30a & vbd & v30e & v29f & v30f & v310;
wire rnx2x7 = rnx2x6 || v311;
wire onx2x7 = onx2x6 || ( rnx2x6 && v311);
wire [7:0] v312 = instruction_bits[31: 24];
wire [7:0] pad_787 = (v312[7:7] == 1'b1) ?24'b111111111111111111111111 : 24'b000000000000000000000000;
wire [31:0] v313 = { pad_787, v312 };
wire v315 = v313 == Advice_4;
wire v316 = v2f0 == Advice_3;
wire [2:0] v317 = instruction_bits[21: 19];
wire [2:0] v318 = { v317 };
wire v319 = v318 == Advice_6;
wire v31a = v2fc & v2fd & v2fe & v2ff & v300 & v301 & v302 & v303 & v2da & v264 & v267 & v26a & v26d & v270 & v273 & v276 & v2b1 & v27e & v2b2 & v283 & v286 & v289;
wire v31b = v2fa & v31a;
wire v31c = v315 & v306 & v294 & v29f & v316 & v299 & v319 & v31b & vaf & v29d & v30f & v310;
wire rnx2x8 = rnx2x7 || v31c;
wire onx2x8 = onx2x7 || ( rnx2x7 && v31c);
wire [31:0] v31d = 32'b10100000000000000000000000000000;
wire [31:0] v31e = In_register_EIP + v31d;
wire v31f = v31e == Out_register_EIP;
wire v320 = v2fc & v2fd & v2fe & v2ff & v300 & v301 & v302 & v303 & v31f & v264 & v267 & v26a & v26d & v270 & v273 & v276 & v2b1 & v27e & v2b2 & v283 & v286 & v289;
wire v321 = v2fa & v320;
wire [7:0] v322 = instruction_bits[39: 32];
wire [7:0] pad_803 = (v322[7:7] == 1'b1) ?24'b111111111111111111111111 : 24'b000000000000000000000000;
wire [31:0] v323 = { pad_803, v322 };
wire v325 = v323 == Advice_4;
wire [2:0] v326 = instruction_bits[29: 27];
wire [2:0] v327 = { v326 };
wire v328 = v327 == Advice_6;
wire v329 = v2e2 == Advice_3;
wire v32a = v321 & v325 & v306 & v299 & v328 & v294 & vba & v329 & v29d & v29f & v30f & v310;
wire rnx2x9 = rnx2x8 || v32a;
wire onx2x9 = onx2x8 || ( rnx2x8 && v32a);
wire [15:0] v32b = instruction_bits[39: 24];
wire [15:0] pad_812 = (v32b[15:15] == 1'b1) ?16'b1111111111111111 : 16'b0000000000000000;
wire [31:0] v32c = { pad_812, v32b };
wire v32e = v32c == Advice_4;
wire [31:0] v330 = ( Advice_13 == 3'd0) ? In_register_EAX :
	( Advice_13 == 3'd1) ? In_register_ECX :
	( Advice_13 == 3'd2) ? In_register_EDX :
	( Advice_13 == 3'd3) ? In_register_EBX :
	( Advice_13 == 3'd4) ? In_register_ESP :
	( Advice_13 == 3'd5) ? In_register_EBP :
	( Advice_13 == 3'd6) ? In_register_ESI : In_register_EDI;
wire [15:0] v331 = v330[31: 16];
wire [31:0] v332 = { v331 , v23e };
wire v333 = v332 == v2f9;
wire v334 = v2fc & v2fd & v2fe & v2ff & v300 & v301 & v302 & v303 & v31f & v264 & v267 & v26a & v26d & v270 & v273 & v276 & v27b & v27e & v280 & v283 & v286 & v289;
wire v335 = v333 & v334;
wire v336 = v2df == Advice_10;
wire v337 = Advice_6 == Advice_13;
wire v338 = v32e & v299 & v335 & v336 & v294 & v316 & v319 & va6 & v29d & v29f & v30f & v310 & v337;
wire rnx2x10 = rnx2x9 || v338;
wire onx2x10 = onx2x9 || ( rnx2x9 && v338);
wire v339 = v2fc & v2fd & v2fe & v2ff & v300 & v301 & v302 & v303 & v2ac & v264 & v267 & v26a & v26d & v270 & v273 & v276 & v27b & v27e & v280 & v283 & v286 & v289;
wire v33a = v333 & v339;
wire [15:0] v33b = instruction_bits[47: 32];
wire [15:0] pad_828 = (v33b[15:15] == 1'b1) ?16'b1111111111111111 : 16'b0000000000000000;
wire [31:0] v33c = { pad_828, v33b };
wire v33e = v33c == Advice_4;
wire v33f = v33a & v33e & v336 & v299 & v29d & v329 & v29f & v328 & v294 & v68 & v30f & v310 & v337;
wire rnx2x11 = rnx2x10 || v33f;
wire onx2x11 = onx2x10 || ( rnx2x10 && v33f);
wire v340 = v2fc & v2fd & v2fe & v2ff & v300 & v301 & v302 & v303 & v2ac & v264 & v267 & v26a & v26d & v270 & v273 & v276 & v2b1 & v27e & v2b2 & v283 & v286 & v289;
wire v341 = v2fa & v340;
wire v342 = v2a1 == Advice_4;
wire v343 = v341 & v342 & v294 & v299 & v29f & v307 & v30a & vb4 & v306 & v29d & v30f & v310;
wire rnx2x12 = rnx2x11 || v343;
wire onx2x12 = onx2x11 || ( rnx2x11 && v343);
wire v344 = v2bb == Advice_4;
wire v345 = v2fc & v2fd & v2fe & v2ff & v300 & v301 & v302 & v303 & v2b9 & v264 & v267 & v26a & v26d & v270 & v273 & v276 & v2b1 & v27e & v2b2 & v283 & v286 & v289;
wire v346 = v2fa & v345;
wire v347 = v344 & v306 & v346 & v319 & v316 & v294 & v299 & v29f & vb7 & v29d & v30f & v310;
wire rnx2x13 = rnx2x12 || v347;
wire onx2x13 = onx2x12 || ( rnx2x12 && v347);
wire v348 = v28f == Advice_4;
wire v349 = v2fc & v2fd & v2fe & v2ff & v300 & v301 & v302 & v303 & v261 & v264 & v267 & v26a & v26d & v270 & v273 & v276 & v2b1 & v27e & v2b2 & v283 & v286 & v289;
wire v34a = v2fa & v349;
wire v34b = v348 & v306 & v294 & v299 & v34a & v29f & v329 & v328 & vac & v29d & v30f & v310;
wire rnx2x14 = rnx2x13 || v34b;
wire onx2x14 = onx2x13 || ( rnx2x13 && v34b);
wire v34c =  v2b4 == memory_0[15: 12] && Advice_10 == memory_0[79: 16] && In_timestamp == memory_0[207: 144] && 4'd0 == memory_0[11: 8] && 1'b1 == memory_0[0: 0] && 6'b000000 == memory_0[7: 2] && 1'b0 == memory_0[1: 1];
wire v34d = v2ec == Advice_7;
wire [31:0] v34f = ( Advice_14 == 3'd0) ? In_register_DSBASE :
	( Advice_14 == 3'd1) ? In_register_DSBASE :
	( Advice_14 == 3'd2) ? In_register_DSBASE :
	( Advice_14 == 3'd3) ? In_register_DSBASE :
	( Advice_14 == 3'd4) ? In_register_SSBASE :
	( Advice_14 == 3'd5) ? In_register_SSBASE :
	( Advice_14 == 3'd6) ? In_register_DSBASE : In_register_DSBASE;
wire [31:0] v350 = v34f + v2dd;
wire [31:0] v351 = v350 + v28d;
wire [31:0] v352 = v351 + v128;
wire v353 = v352 == Advice_10;
wire v354 = Advice_7 == Advice_14;
wire v355 = v299 & v34c & v34d & v294 & v307 & v30a & v30e & v1aa & v353 & v29d & v305 & v29f & v30f & v354 & v310;
wire rnx2x15 = rnx2x14 || v355;
wire onx2x15 = onx2x14 || ( rnx2x14 && v355);
wire [31:0] v356 = v351 + v30c;
wire v357 = v356 == Advice_10;
wire v358 = v31b & v299 & v102 & v34d & v357 & v307 & v315 & v294 & v30a & v34c & v29d & v29f & v30f & v354 & v310;
wire rnx2x16 = rnx2x15 || v358;
wire onx2x16 = onx2x15 || ( rnx2x15 && v358);
wire [7:0] v359 = instruction_bits[55: 48];
wire [7:0] pad_858 = (v359[7:7] == 1'b1) ?24'b111111111111111111111111 : 24'b000000000000000000000000;
wire [31:0] v35a = { pad_858, v359 };
wire v35c = v35a == Advice_4;
wire [31:0] v35d = v351 + v2a1;
wire v35e = v35d == Advice_10;
wire v35f = v346 & v35c & v294 & v299 & v30a & v34c & v35e & v34d & v307 & v29f & v124 & v29d & v30f & v354 & v310;
wire rnx2x17 = rnx2x16 || v35f;
wire onx2x17 = onx2x16 || ( rnx2x16 && v35f);
wire v360 = v2a3 == Advice_10;
wire v361 = v35c & v360 & v294 & v29d & v34c & v299 & v30a & v346 & v141 & v29f & v310;
wire rnx2x18 = rnx2x17 || v361;
wire onx2x18 = onx2x17 || ( rnx2x17 && v361);
wire v362 = v2f0 == Advice_7;
wire [31:0] v363 = { 30'b000000000000000000000000000000, va1 };
wire [31:0] v365 = v330 << v363;
wire [31:0] v366 = v350 + v365;
wire [31:0] v367 = v366 + v128;
wire v368 = v367 == Advice_10;
wire v369 = v318 == Advice_2;
wire v36a = Advice_2 == Advice_13;
wire v36b = v31b & v315 & v34c & v15e & v362 & v368 & v369 & v30a & v299 & v316 & v29f & v294 & v29d & v30f & v36a & v354 & v310;
wire rnx2x19 = rnx2x18 || v36b;
wire onx2x19 = onx2x18 || ( rnx2x18 && v36b);
wire [7:0] v36c = instruction_bits[63: 56];
wire [7:0] pad_877 = (v36c[7:7] == 1'b1) ?24'b111111111111111111111111 : 24'b000000000000000000000000;
wire [31:0] v36d = { pad_877, v36c };
wire v36f = v36d == Advice_4;
wire [31:0] v370 = v366 + v2bb;
wire v371 = v370 == Advice_10;
wire v372 = v34a & v36f & v294 & v34c & v299 & v371 & v362 & v369 & v29f & v316 & v171 & v30a & v29d & v30f & v36a & v354 & v310;
wire rnx2x20 = rnx2x19 || v372;
wire onx2x20 = onx2x19 || ( rnx2x19 && v372);
wire [31:0] v373 = v366 + v313;
wire v374 = v373 == Advice_10;
wire v375 = v374 & v325 & v299 & v294 & v34c & v369 & v316 & v29f & v321 & v30a & v362 & v174 & v29d & v30f & v36a & v354 & v310;
wire rnx2x21 = rnx2x20 || v375;
wire onx2x21 = onx2x20 || ( rnx2x20 && v375);
wire [31:0] v377 = ( Advice_15 == 2'd0) ? In_register_EDX :
	( Advice_15 == 2'd1) ? In_register_ESI :
	( Advice_15 == 2'd2) ? In_register_EBX : In_register_EDI;
wire [31:0] v378 = v377 << v363;
wire [31:0] v379 = v28c + v378;
wire [31:0] v37a = v379 + v2bb;
wire v37b = v37a == Advice_10;
wire v37d = instruction_bits[19: 19];
wire v37c = instruction_bits[21: 21];
wire [1:0] v37e = { v37d , v37c };
wire v380 = v37e == Advice_16;
wire v381 = Advice_16 == Advice_15;
wire v382 = v34a & v36f & v37b & v294 & v299 & v34c & v29d & v380 & v121 & v30a & v29f & v381 & v310;
wire rnx2x22 = rnx2x21 || v382;
wire onx2x22 = onx2x21 || ( rnx2x21 && v382);
wire [31:0] v383 = v351 + v2bb;
wire v384 = v383 == Advice_10;
wire v385 = v34a & v183 & v36f & v294 & v299 & v34c & v362 & v316 & v30a & v29d & v384 & v29f & v30f & v354 & v310;
wire rnx2x23 = rnx2x22 || v385;
wire onx2x23 = onx2x22 || ( rnx2x22 && v385);
wire v386 = v31b & v362 & v353 & v34c & v294 & v29f & v30a & v315 & v316 & v185 & v299 & v29d & v30f & v354 & v310;
wire rnx2x24 = rnx2x23 || v386;
wire onx2x24 = onx2x23 || ( rnx2x23 && v386);
wire [31:0] v387 = v351 + v313;
wire v388 = v387 == Advice_10;
wire v389 = v294 & v325 & v299 & v29f & v34c & v316 & v30a & v187 & v321 & v388 & v29d & v362 & v30f & v354 & v310;
wire rnx2x25 = rnx2x24 || v389;
wire onx2x25 = onx2x24 || ( rnx2x24 && v389);
wire [31:0] v38b = ( Advice_17 == 3'd0) ? In_register_ESBASE :
	( Advice_17 == 3'd1) ? In_register_ESBASE :
	( Advice_17 == 3'd2) ? In_register_ESBASE :
	( Advice_17 == 3'd3) ? In_register_ESBASE :
	( Advice_17 == 3'd4) ? In_register_ESBASE :
	( Advice_17 == 3'd5) ? In_register_ESBASE :
	( Advice_17 == 3'd6) ? In_register_ESBASE : In_register_ESBASE;
wire [31:0] v38c = v38b + v2dd;
wire [31:0] v38d = v38c + v28d;
wire [31:0] v38e = v38d + v2bb;
wire v38f = v38e == Advice_10;
wire v390 = Advice_7 == Advice_17;
wire v391 = v34a & v319 & v36f & v38f & v299 & v34c & v362 & v29f & v1a8 & v316 & v294 & v29d & v30f & v390 & v310;
wire rnx2x26 = rnx2x25 || v391;
wire onx2x26 = onx2x25 || ( rnx2x25 && v391);
wire [31:0] v393 = ( Advice_18 == 3'd0) ? In_register_EBX :
	( Advice_18 == 3'd1) ? In_register_EBX :
	( Advice_18 == 3'd2) ? In_register_EBP :
	( Advice_18 == 3'd3) ? In_register_EBP :
	( Advice_18 == 3'd4) ? In_register_ESI :
	( Advice_18 == 3'd5) ? In_register_EDI :
	( Advice_18 == 3'd6) ? In_register_EBP : In_register_EBX;
wire [31:0] v394 = v393 & v2de;
wire [31:0] v395 = v34f + v394;
wire [31:0] v397 = ( Advice_19 == 1'd0) ? In_register_ESI : In_register_EDI;
wire [31:0] v398 = v397 & v2de;
wire [31:0] v399 = 32'b10000000000000000000000000000000;
wire [31:0] v39b = v398 << v399;
wire [31:0] v39c = v395 + v39b;
wire [31:0] v39d = v39c + v32c;
wire [15:0] v39e = v39d[15:0];
wire [31:0] v39f = { 16'b0000000000000000, v39e };
wire v3a0 = v39f == Advice_10;
wire v3a1 = { v57 };
wire v3a3 = v3a1 == Advice_20;
wire [7:0] v3a4 = instruction_bits[47: 40];
wire [7:0] pad_933 = (v3a4[7:7] == 1'b1) ?24'b111111111111111111111111 : 24'b000000000000000000000000;
wire [31:0] v3a5 = { pad_933, v3a4 };
wire v3a7 = v3a5 == Advice_4;
wire v3a8 = v3a1 == Advice_8;
wire v3a9 = instruction_bits[16: 16];
wire v3aa = { v3a9 };
wire v3ac = v3aa == Advice_21;
wire [2:0] v3ad = { Advice_8 , vd8 };
wire v3ae = v3ad == Advice_18;
wire v3af = Advice_21 == Advice_19;
wire [2:0] v3b0 = { Advice_20 , vd8 };
wire v3b1 = v3b0 == Advice_14;
wire v3b2 = v341 & v3a0 & v299 & v34c & v29d & v3a3 & v29f & v294 & v11c & v319 & v3a7 & v3a8 & v3ac & v3ae & v3af & v3b1 & v310;
wire rnx2x27 = rnx2x26 || v3b2;
wire onx2x27 = onx2x26 || ( rnx2x26 && v3b2);
wire [7:0] v3b3 = instruction_bits[71: 64];
wire [7:0] pad_948 = (v3b3[7:7] == 1'b1) ?24'b111111111111111111111111 : 24'b000000000000000000000000;
wire [31:0] v3b4 = { pad_948, v3b3 };
wire v3b6 = v3b4 == Advice_4;
wire [31:0] v3b7 = { 30'b000000000000000000000000000000, v66 };
wire [31:0] v3b9 = v330 << v3b7;
wire [31:0] v3ba = v38c + v3b9;
wire [31:0] v3bb = v3ba + v28f;
wire v3bc = v3bb == Advice_10;
wire v3bd = v327 == Advice_2;
wire v3be = v2e2 == Advice_7;
wire [31:0] v3bf = 32'b10010000000000000000000000000000;
wire [31:0] v3c0 = In_register_EIP + v3bf;
wire v3c1 = v3c0 == Out_register_EIP;
wire v3c2 = v2fc & v2fd & v2fe & v2ff & v300 & v301 & v302 & v303 & v3c1 & v264 & v267 & v26a & v26d & v270 & v273 & v276 & v2b1 & v27e & v2b2 & v283 & v286 & v289;
wire v3c3 = v2fa & v3c2;
wire v3c4 = v3b6 & v319 & v34c & v3bc & v3bd & v3be & v294 & v329 & v152 & v29d & v299 & v3c3 & v29f & v30f & v36a & v390 & v310;
wire rnx2x28 = rnx2x27 || v3c4;
wire onx2x28 = onx2x27 || ( rnx2x27 && v3c4);
wire v3c5 = v2bd == Advice_10;
wire v3c6 = v34a & v3c5 & v294 & v36f & v34c & v30a & v18a & v299 & v29d & v29f & v310;
wire rnx2x29 = rnx2x28 || v3c6;
wire onx2x29 = onx2x28 || ( rnx2x28 && v3c6);
wire [31:0] v3c7 = In_register_FSBASE + v128;
wire [31:0] v3c8 = v3c7 + v28d;
wire [31:0] v3c9 = v3c8 + v2bb;
wire v3ca = v3c9 == Advice_10;
wire v3cb = v34a & v3ca & v294 & v299 & v34c & v319 & v1a7 & v36f & v29d & v29f & v310;
wire rnx2x30 = rnx2x29 || v3cb;
wire onx2x30 = onx2x29 || ( rnx2x29 && v3cb);
wire [31:0] v3cc = v38b + v377;
wire [31:0] v3cd = v3cc + v28d;
wire [31:0] v3ce = v3cd + v128;
wire v3cf = v3ce == Advice_10;
wire [1:0] v3d0 = { v3a9 , v114 };
wire v3d2 = v3d0 == Advice_22;
wire v3d4 = v3d0 == Advice_23;
wire v3d5 = Advice_23 == Advice_15;
wire [2:0] v3d6 = { Advice_22 , v11 };
wire v3d7 = v3d6 == Advice_17;
wire v3d8 = v31b & v299 & v34c & v315 & v3cf & v3d2 & v29f & v294 & v3d4 & v319 & v14c & v29d & v3d5 & v3d7 & v310;
wire rnx2x31 = rnx2x30 || v3d8;
wire onx2x31 = onx2x30 || ( rnx2x30 && v3d8);
wire [31:0] v3d9 = v38d + v313;
wire v3da = v3d9 == Advice_10;
wire v3db = v294 & v299 & v34c & v362 & v29f & v100 & v316 & v321 & v319 & v3da & v325 & v29d & v30f & v390 & v310;
wire rnx2x32 = rnx2x31 || v3db;
wire onx2x32 = onx2x31 || ( rnx2x31 && v3db);
wire [31:0] v3dd = ( Advice_24 == 3'd0) ? In_register_FSBASE :
	( Advice_24 == 3'd1) ? In_register_FSBASE :
	( Advice_24 == 3'd2) ? In_register_FSBASE :
	( Advice_24 == 3'd3) ? In_register_FSBASE :
	( Advice_24 == 3'd4) ? In_register_FSBASE :
	( Advice_24 == 3'd5) ? In_register_FSBASE :
	( Advice_24 == 3'd6) ? In_register_FSBASE : In_register_FSBASE;
wire [31:0] v3de = v3dd + v2dd;
wire [31:0] v3df = v3de + v3b9;
wire [31:0] v3e0 = v3df + v323;
wire v3e1 = v3e0 == Advice_10;
wire v3e2 = Advice_7 == Advice_24;
wire v3e3 = v341 & v3a7 & v29d & v3be & v3e1 & v299 & v294 & v319 & v34c & v17e & v329 & v3bd & v29f & v30f & v36a & v3e2 & v310;
wire rnx2x33 = rnx2x32 || v3e3;
wire onx2x33 = onx2x32 || ( rnx2x32 && v3e3);
wire [31:0] v3e5 = ( Advice_25 == 2'd0) ? In_register_DSBASE :
	( Advice_25 == 2'd1) ? In_register_DSBASE :
	( Advice_25 == 2'd2) ? In_register_DSBASE : In_register_DSBASE;
wire [31:0] v3e7 = ( Advice_26 == 1'd0) ? In_register_EDI : In_register_EBX;
wire [31:0] v3e8 = v3e7 & v2de;
wire [31:0] v3e9 = v3e5 + v3e8;
wire [31:0] v3ea = v3e9 + v28d;
wire [31:0] v3eb = v3ea + v128;
wire [15:0] v3ec = v3eb[15:0];
wire [31:0] v3ed = { 16'b0000000000000000, v3ec };
wire v3ee = v3ed == Advice_10;
wire v3ef = Advice_8 == Advice_26;
wire [1:0] v3f0 = { Advice_20 , v11 };
wire v3f1 = v3f0 == Advice_25;
wire v3f2 = v31b & v3ee & v315 & v294 & v3a3 & v178 & v3a8 & v34c & v319 & v29d & v299 & v29f & v3ef & v3f1 & v310;
wire rnx2x34 = rnx2x33 || v3f2;
wire onx2x34 = onx2x33 || ( rnx2x33 && v3f2);
wire [31:0] v3f3 = v39c + v313;
wire [15:0] v3f4 = v3f3[15:0];
wire [31:0] v3f5 = { 16'b0000000000000000, v3f4 };
wire v3f6 = v3f5 == Advice_10;
wire v3f7 = v321 & v325 & v294 & v29d & v299 & v3a3 & v3ac & v319 & v3f6 & v3a8 & v186 & v34c & v29f & v3ae & v3af & v3b1 & v310;
wire rnx2x35 = rnx2x34 || v3f7;
wire onx2x35 = onx2x34 || ( rnx2x34 && v3f7);
wire [31:0] v3f8 = v39c + v128;
wire [15:0] v3f9 = v3f8[15:0];
wire [31:0] v3fa = { 16'b0000000000000000, v3f9 };
wire v3fb = v3fa == Advice_10;
wire v3fc = v31b & v315 & v3a3 & v3ac & v142 & v3fb & v3a8 & v29f & v319 & v294 & v299 & v34c & v29d & v3ae & v3af & v3b1 & v310;
wire rnx2x36 = rnx2x35 || v3fc;
wire onx2x36 = onx2x35 || ( rnx2x35 && v3fc);
wire [15:0] v3fd = 16'b0000000111111111;
wire [15:0] v3fe = v2c2 + v3fd;
wire [15:0] v3ff = 16'b0000000011111111;
wire v400 = v3fe < v3ff;
wire v401 = v400 == Out_register_CF;
wire v402 = v400 == Out_register_OF;
wire v403 = v2ce & v245 & v248 & v2cf & v253 & v256 & v259 & v25c & v2b9 & v264 & v267 & v26a & v26d & v270 & v273 & v276 & v401 & v27e & v402 & v283 & v286 & v289;
wire v404 = v370 == Advice_5;
wire v405 = v2f0 == Advice_2;
wire v406 = v318 == Advice_3;
wire v407 = Advice_3 == Advice_13;
wire v408 = Advice_2 == Advice_14;
wire v409 = v403 & v404 & v2d6 & v405 & v299 & v406 & v294 & v2f1 & v8e & v29d & v29f & v2e4 & v407 & v408;
wire rnx2x37 = rnx2x36 || v409;
wire onx2x37 = onx2x36 || ( rnx2x36 && v409);
wire v40b = instruction_bits[24: 24];
wire v40a = instruction_bits[26: 26];
wire [1:0] v40c = { v40b , v40a };
wire v40d = v40c == Advice_22;
wire v40e = v40c == Advice_23;
wire [31:0] v40f = v2dd << v3b7;
wire [31:0] v410 = v3cc + v40f;
wire [31:0] v411 = v410 + v128;
wire v412 = v411 == Advice_10;
wire v413 = Advice_2 == Advice_11;
wire v414 = v321 & v325 & v299 & v319 & v294 & v34c & v40d & v3bd & v29f & v40e & v412 & v190 & v29d & v3d5 & v413 & v3d7 & v310;
wire rnx2x38 = rnx2x37 || v414;
wire onx2x38 = onx2x37 || ( rnx2x37 && v414);
wire v415 =  v295 == memory_0[15: 12] && Advice_10 == memory_0[79: 16] && In_timestamp == memory_0[207: 144] && 4'd0 == memory_0[11: 8] && 1'b1 == memory_0[0: 0] && 6'b000000 == memory_0[7: 2] && 1'b0 == memory_0[1: 1];
wire [15:0] v416 = instruction_bits[71: 56];
wire [15:0] pad_1047 = (v416[15:15] == 1'b1) ?16'b1111111111111111 : 16'b0000000000000000;
wire [31:0] v417 = { pad_1047, v416 };
wire v419 = v417 == Advice_4;
wire v41a = v2fc & v2fd & v2fe & v2ff & v300 & v301 & v302 & v303 & v3c1 & v264 & v267 & v26a & v26d & v270 & v273 & v276 & v27b & v27e & v280 & v283 & v286 & v289;
wire v41b = v333 & v41a;
wire v41c = v384 & v299 & v29f & v415 & v419 & v294 & v362 & v316 & v41b & v29d & v319 & v1f3 & v30f & v354 & v310 & v337;
wire rnx2x39 = rnx2x38 || v41c;
wire onx2x39 = onx2x38 || ( rnx2x38 && v41c);
wire [15:0] v41d = instruction_bits[79: 64];
wire [15:0] pad_1054 = (v41d[15:15] == 1'b1) ?16'b1111111111111111 : 16'b0000000000000000;
wire [31:0] v41e = { pad_1054, v41d };
wire v420 = v41e == Advice_4;
wire [31:0] v422 = ( Advice_27 == 3'd0) ? In_register_EAX :
	( Advice_27 == 3'd1) ? In_register_ECX :
	( Advice_27 == 3'd2) ? In_register_EDX :
	( Advice_27 == 3'd3) ? In_register_EBX :
	( Advice_27 == 3'd4) ? In_register_ESP :
	( Advice_27 == 3'd5) ? In_register_EBP :
	( Advice_27 == 3'd6) ? In_register_ESI : In_register_EDI;
wire [15:0] v423 = v422[31: 16];
wire [31:0] v424 = { v423 , v23e };
wire v425 = v424 == v2f9;
wire [31:0] v426 = 32'b01010000000000000000000000000000;
wire [31:0] v427 = In_register_EIP + v426;
wire v428 = v427 == Out_register_EIP;
wire v429 = v2fc & v2fd & v2fe & v2ff & v300 & v301 & v302 & v303 & v428 & v264 & v267 & v26a & v26d & v270 & v273 & v276 & v27b & v27e & v280 & v283 & v286 & v289;
wire v42a = v425 & v429;
wire [31:0] v42b = v350 + v3b9;
wire [31:0] v42c = v42b + v28f;
wire v42d = v42c == Advice_10;
wire v42e = Advice_6 == Advice_27;
wire v42f = v420 & v42a & v415 & v42d & v299 & v3bd & v329 & v319 & v1b5 & v29f & v294 & v29d & v3be & v30f & v36a & v354 & v310 & v42e;
wire rnx2x40 = rnx2x39 || v42f;
wire onx2x40 = onx2x39 || ( rnx2x39 && v42f);
wire [31:0] v430 = v3e5 + v377;
wire [31:0] v431 = v430 + v28d;
wire [31:0] v432 = v431 + v128;
wire v433 = v432 == Advice_10;
wire [15:0] v434 = v2dd[31: 16];
wire [31:0] v435 = { v434 , v23e };
wire v436 = v435 == v2f9;
wire v437 = v436 & v334;
wire v438 = Advice_22 == Advice_25;
wire v439 = v299 & v32e & v294 & v433 & v415 & v29f & vdb & v3d4 & v437 & v319 & v3d2 & v29d & v3d5 & v438 & v310 & v2e4;
wire rnx2x41 = rnx2x40 || v439;
wire onx2x41 = onx2x40 || ( rnx2x40 && v439);
wire v43a = v388 & v316 & v294 & v33a & v299 & v33e & v415 & v205 & v319 & v362 & v29d & v29f & v30f & v354 & v310 & v337;
wire rnx2x42 = rnx2x41 || v43a;
wire onx2x42 = onx2x41 || ( rnx2x41 && v43a);
wire v43b = v2fc & v2fd & v2fe & v2ff & v300 & v301 & v302 & v303 & v2b9 & v264 & v267 & v26a & v26d & v270 & v273 & v276 & v27b & v27e & v280 & v283 & v286 & v289;
wire v43c = v425 & v43b;
wire [15:0] v43d = instruction_bits[55: 40];
wire [15:0] pad_1086 = (v43d[15:15] == 1'b1) ?16'b1111111111111111 : 16'b0000000000000000;
wire [31:0] v43e = { pad_1086, v43d };
wire v440 = v43e == Advice_4;
wire [31:0] v441 = v42b + v323;
wire v442 = v441 == Advice_10;
wire v443 = v43c & v440 & v29d & v415 & v3bd & v3be & v329 & v319 & v1b1 & v299 & v442 & v294 & v29f & v30f & v36a & v354 & v310 & v42e;
wire rnx2x43 = rnx2x42 || v443;
wire onx2x43 = onx2x42 || ( rnx2x42 && v443);
wire v444 = v33e & v33a & v294 & v29f & v299 & v415 & v3be & v319 & v329 & v353 & v1dc & v29d & v30f & v354 & v310 & v337;
wire rnx2x44 = rnx2x43 || v444;
wire onx2x44 = onx2x43 || ( rnx2x43 && v444);
wire v445 = v2fc & v2fd & v2fe & v2ff & v300 & v301 & v302 & v303 & v428 & v264 & v267 & v26a & v26d & v270 & v273 & v276 & v2b1 & v27e & v2b2 & v283 & v286 & v289;
wire v446 = v2fa & v445;
wire [31:0] v447 = instruction_bits[79: 48];
wire v449 = v447 == Advice_4;
wire v44b = instruction_bits[8: 8];
wire v44a = instruction_bits[10: 10];
wire [1:0] v44c = { v44b , v44a };
wire v44d = v44c == Advice_22;
wire v44e = v44c == Advice_23;
wire [31:0] v44f = v431 + v2a1;
wire v450 = v44f == Advice_10;
wire v451 = v446 & v449 & v294 & v299 & v44d & v30a & v44e & v135 & v29d & v450 & v34c & v29f & v3d5 & v438 & v310;
wire rnx2x45 = rnx2x44 || v451;
wire onx2x45 = onx2x44 || ( rnx2x44 && v451);
wire v452 = v341 & v294 & v342 & v353 & v34d & v299 & v34c & v307 & v29f & v30a & v172 & v29d & v30f & v354 & v310;
wire rnx2x46 = rnx2x45 || v452;
wire onx2x46 = onx2x45 || ( rnx2x45 && v452);
wire v453 = v446 & v360 & v34c & v299 & v111 & v449 & v30a & v294 & v29d & v29f & v310;
wire rnx2x47 = rnx2x46 || v453;
wire onx2x47 = onx2x46 || ( rnx2x46 && v453);
wire v454 = v346 & v344 & v29d & v299 & v34c & v34d & v294 & v307 & v30a & v357 & v134 & v29f & v30f & v354 & v310;
wire rnx2x48 = rnx2x47 || v454;
wire onx2x48 = onx2x47 || ( rnx2x47 && v454);
wire v455 = v346 & v30a & v368 & v299 & v362 & v369 & v34c & v10b & v316 & v29d & v344 & v294 & v29f & v30f & v36a & v354 & v310;
wire rnx2x49 = rnx2x48 || v455;
wire onx2x49 = onx2x48 || ( rnx2x48 && v455);
wire v456 = v348 & v374 & v294 & v29f & v299 & v34c & v34a & v14e & v362 & v369 & v30a & v316 & v29d & v30f & v36a & v354 & v310;
wire rnx2x50 = rnx2x49 || v456;
wire onx2x50 = onx2x49 || ( rnx2x49 && v456);
wire [31:0] v457 = instruction_bits[87: 56];
wire v459 = v457 == Advice_4;
wire [31:0] v45a = 32'b11010000000000000000000000000000;
wire [31:0] v45b = In_register_EIP + v45a;
wire v45c = v45b == Out_register_EIP;
wire v45d = v2fc & v2fd & v2fe & v2ff & v300 & v301 & v302 & v303 & v45c & v264 & v267 & v26a & v26d & v270 & v273 & v276 & v2b1 & v27e & v2b2 & v283 & v286 & v289;
wire v45e = v2fa & v45d;
wire v45f = v459 & v371 & v294 & v299 & v34c & v369 & v362 & v45e & v17f & v316 & v30a & v29d & v29f & v30f & v36a & v354 & v310;
wire rnx2x51 = rnx2x50 || v45f;
wire onx2x51 = onx2x50 || ( rnx2x50 && v45f);
wire v460 = v45e & v362 & v30a & v34c & v384 & v316 & v29d & v299 & v13e & v459 & v294 & v29f & v30f & v354 & v310;
wire rnx2x52 = rnx2x51 || v460;
wire onx2x52 = onx2x51 || ( rnx2x51 && v460);
wire v461 = v299 & v362 & v344 & v1a9 & v316 & v346 & v353 & v30a & v294 & v34c & v29d & v29f & v30f & v354 & v310;
wire rnx2x53 = rnx2x52 || v461;
wire onx2x53 = onx2x52 || ( rnx2x52 && v461);
wire v462 = v34a & v348 & v388 & v294 & v362 & v299 & v316 & v29f & v30a & v34c & v153 & v29d & v30f & v354 & v310;
wire rnx2x54 = rnx2x53 || v462;
wire onx2x54 = onx2x53 || ( rnx2x53 && v462);
wire [31:0] v463 = v2dd << v363;
wire [31:0] v464 = v28c + v463;
wire [31:0] v465 = v464 + v2bb;
wire v466 = v465 == Advice_10;
wire v467 = v299 & v294 & v34c & v173 & v369 & v459 & v30a & v45e & v466 & v29d & v29f & v413 & v310;
wire rnx2x55 = rnx2x54 || v467;
wire onx2x55 = onx2x54 || ( rnx2x54 && v467);
wire [31:0] v469 = ( Advice_28 == 3'd0) ? In_register_DSBASE :
	( Advice_28 == 3'd1) ? In_register_DSBASE :
	( Advice_28 == 3'd2) ? In_register_SSBASE :
	( Advice_28 == 3'd3) ? In_register_SSBASE :
	( Advice_28 == 3'd4) ? In_register_DSBASE :
	( Advice_28 == 3'd5) ? In_register_DSBASE :
	( Advice_28 == 3'd6) ? In_register_SSBASE : In_register_DSBASE;
wire [31:0] v46a = v469 + v394;
wire [31:0] v46c = ( Advice_29 == 3'd0) ? In_register_ESI :
	( Advice_29 == 3'd1) ? In_register_EDI :
	( Advice_29 == 3'd2) ? In_register_ESI :
	( Advice_29 == 3'd3) ? In_register_EDI :
	( Advice_29 == 3'd4) ? v128 :
	( Advice_29 == 3'd5) ? v128 :
	( Advice_29 == 3'd6) ? v128 : v128;
wire [31:0] v46d = v46c & v2de;
wire [31:0] v46e = v46d << v399;
wire [31:0] v46f = v46a + v46e;
wire [31:0] v470 = v46f + v32c;
wire [15:0] v471 = v470[15:0];
wire [31:0] v472 = { 16'b0000000000000000, v471 };
wire v473 = v472 == Advice_10;
wire [31:0] v474 = instruction_bits[71: 40];
wire v476 = v474 == Advice_4;
wire v477 = Advice_3 == Advice_18;
wire v478 = Advice_2 == Advice_29;
wire v479 = Advice_7 == Advice_28;
wire v47a = v3c3 & v473 & v316 & v299 & v362 & v34c & v319 & v405 & v29d & v294 & v476 & v12f & v29f & v477 & v478 & v479 & v310;
wire rnx2x56 = rnx2x55 || v47a;
wire onx2x56 = onx2x55 || ( rnx2x55 && v47a);
wire v47b = v45e & v294 & v299 & v459 & v362 & v38f & v34c & v319 & v29d & v182 & v316 & v29f & v30f & v390 & v310;
wire rnx2x57 = rnx2x56 || v47b;
wire onx2x57 = onx2x56 || ( rnx2x56 && v47b);
wire [31:0] v47c = v3de + v28d;
wire [31:0] v47d = v47c + v128;
wire v47e = v47d == Advice_10;
wire v47f = v346 & v299 & v362 & v34c & v344 & v47e & v294 & v29d & v319 & v316 & v19a & v29f & v30f & v3e2 & v310;
wire rnx2x58 = rnx2x57 || v47f;
wire onx2x58 = onx2x57 || ( rnx2x57 && v47f);
wire [31:0] v481 = ( Advice_30 == 3'd0) ? In_register_GSBASE :
	( Advice_30 == 3'd1) ? In_register_GSBASE :
	( Advice_30 == 3'd2) ? In_register_GSBASE :
	( Advice_30 == 3'd3) ? In_register_GSBASE :
	( Advice_30 == 3'd4) ? In_register_GSBASE :
	( Advice_30 == 3'd5) ? In_register_GSBASE :
	( Advice_30 == 3'd6) ? In_register_GSBASE : In_register_GSBASE;
wire [31:0] v482 = v481 + v2dd;
wire [31:0] v483 = v377 << v3b7;
wire [31:0] v484 = v482 + v483;
wire [31:0] v485 = v484 + v323;
wire v486 = v485 == Advice_10;
wire v488 = instruction_bits[27: 27];
wire v487 = instruction_bits[29: 29];
wire [1:0] v489 = { v488 , v487 };
wire v48a = v489 == Advice_16;
wire v48b = Advice_7 == Advice_30;
wire v48c = v3c3 & v476 & v486 & v299 & v3be & v48a & v34c & v319 & v29d & v15d & v294 & v329 & v29f & v30f & v381 & v48b & v310;
wire rnx2x59 = rnx2x58 || v48c;
wire onx2x59 = onx2x58 || ( rnx2x58 && v48c);
wire v48d = v3c5 & v294 & v299 & v30a & v29f & v12b & v459 & v34c & v45e & v29d & v310;
wire rnx2x60 = rnx2x59 || v48d;
wire onx2x60 = onx2x59 || ( rnx2x59 && v48d);
wire [31:0] v48e = v3dd + v377;
wire [31:0] v48f = v48e + v28d;
wire [31:0] v490 = v48f + v313;
wire v491 = v490 == Advice_10;
wire v492 = v3d6 == Advice_24;
wire v493 = v34a & v34c & v299 & v348 & v491 & v294 & v3d4 & v29f & v319 & v3d2 & v17b & v29d & v3d5 & v492 & v310;
wire rnx2x61 = rnx2x60 || v493;
wire onx2x61 = onx2x60 || ( rnx2x60 && v493);
wire v494 = v346 & v34c & v3ee & v299 & v319 & v3a3 & v3a8 & v344 & v294 & v199 & v29d & v29f & v3ef & v3f1 & v310;
wire rnx2x62 = rnx2x61 || v494;
wire onx2x62 = onx2x61 || ( rnx2x61 && v494);
wire [31:0] v495 = v46f + v313;
wire [15:0] v496 = v495[15:0];
wire [31:0] v497 = { 16'b0000000000000000, v496 };
wire v498 = v497 == Advice_10;
wire v499 = v498 & v34a & v299 & v34c & v294 & v405 & v362 & v348 & v316 & v319 & v130 & v29d & v29f & v477 & v478 & v479 & v310;
wire rnx2x63 = rnx2x62 || v499;
wire onx2x63 = onx2x62 || ( rnx2x62 && v499);
wire [31:0] v49a = 32'b00110000000000000000000000000000;
wire [31:0] v49b = In_register_EIP + v49a;
wire v49c = v49b == Out_register_EIP;
wire v49d = v2fc & v2fd & v2fe & v2ff & v300 & v301 & v302 & v303 & v49c & v264 & v267 & v26a & v26d & v270 & v273 & v276 & v2b1 & v27e & v2b2 & v283 & v286 & v289;
wire v49e = v2fa & v49d;
wire [31:0] v4a0 = ( Advice_31 == 3'd0) ? In_register_SSBASE :
	( Advice_31 == 3'd1) ? In_register_SSBASE :
	( Advice_31 == 3'd2) ? In_register_SSBASE :
	( Advice_31 == 3'd3) ? In_register_SSBASE :
	( Advice_31 == 3'd4) ? In_register_SSBASE :
	( Advice_31 == 3'd5) ? In_register_SSBASE :
	( Advice_31 == 3'd6) ? In_register_SSBASE : In_register_SSBASE;
wire [31:0] v4a1 = v4a0 + v2dd;
wire [31:0] v4a2 = v4a1 + v3b9;
wire [31:0] v4a3 = v4a2 + v28f;
wire v4a4 = v4a3 == Advice_10;
wire [31:0] v4a5 = instruction_bits[95: 64];
wire v4a7 = v4a5 == Advice_4;
wire v4a8 = Advice_7 == Advice_31;
wire v4a9 = v49e & v4a4 & v294 & v299 & v34c & v3bd & v196 & v3be & v4a7 & v329 & v319 & v29d & v29f & v30f & v36a & v4a8 & v310;
wire rnx2x64 = rnx2x63 || v4a9;
wire onx2x64 = onx2x63 || ( rnx2x63 && v4a9);
wire [31:0] v4aa = In_register_GSBASE + v128;
wire [31:0] v4ab = v4aa + v28d;
wire [31:0] v4ac = v4ab + v2bb;
wire v4ad = v4ac == Advice_10;
wire v4ae = v45e & v459 & v4ad & v294 & v29d & v161 & v34c & v319 & v299 & v29f & v310;
wire rnx2x65 = rnx2x64 || v4ae;
wire onx2x65 = onx2x64 || ( rnx2x64 && v4ae);
wire [31:0] v4af = v3e5 + v398;
wire [31:0] v4b0 = v4af + v28d;
wire [31:0] v4b1 = v4b0 + v128;
wire [15:0] v4b2 = v4b1[15:0];
wire [31:0] v4b3 = { 16'b0000000000000000, v4b2 };
wire v4b4 = v4b3 == Advice_10;
wire v4b5 = v3aa == Advice_20;
wire v4b6 = v3aa == Advice_8;
wire v4b7 = Advice_8 == Advice_19;
wire v4b8 = v346 & v344 & v4b4 & v294 & v299 & v4b5 & v319 & v34c & v133 & v4b6 & v29d & v29f & v4b7 & v3f1 & v310;
wire rnx2x66 = rnx2x65 || v4b8;
wire onx2x66 = onx2x65 || ( rnx2x65 && v4b8);
wire [31:0] v4b9 = 32'b00000000000000000000000000000000;
wire [31:0] v4ba = ( Advice_1 == 1'd0) ? v4b9 : In_register_EBP;
wire [31:0] v4bb = v4ba & v2de;
wire [31:0] v4bc = v34f + v4bb;
wire [31:0] v4bd = v4bc + v39b;
wire [31:0] v4be = v4bd + v128;
wire [15:0] v4bf = v4be[15:0];
wire [31:0] v4c0 = { 16'b0000000000000000, v4bf };
wire v4c1 = v4c0 == Advice_10;
wire v4c2 = Advice_8 == Advice_1;
wire v4c3 = v344 & v29f & v299 & v346 & v137 & v34c & v3a3 & v3ac & v3a8 & v319 & v294 & v4c1 & v29d & v4c2 & v3af & v3b1 & v310;
wire rnx2x67 = rnx2x66 || v4c3;
wire onx2x67 = onx2x66 || ( rnx2x66 && v4c3);
wire [31:0] v4c4 = v482 + v3b9;
wire [31:0] v4c5 = v4c4 + v128;
wire v4c6 = v4c5 == Advice_10;
wire v4c7 = v34a & v348 & v4c6 & v294 & v3be & v319 & v299 & v3bd & v34c & v329 & v29f & v15a & v29d & v30f & v36a & v48b & v310;
wire rnx2x68 = rnx2x67 || v4c7;
wire onx2x68 = onx2x67 || ( rnx2x67 && v4c7);
wire [31:0] v4c8 = v430 + v463;
wire [31:0] v4c9 = v4c8 + v128;
wire v4ca = v4c9 == Advice_5;
wire v4cb = v3d0 == Advice_16;
wire v4cd = v3d0 == Advice_32;
wire v4ce = v2ce & v245 & v248 & v2cf & v253 & v256 & v259 & v25c & v2f4 & v264 & v267 & v26a & v26d & v270 & v273 & v276 & v401 & v27e & v402 & v283 & v286 & v289;
wire v4cf = Advice_32 == Advice_15;
wire v4d0 = Advice_16 == Advice_25;
wire v4d1 = v299 & v2d6 & v4ca & v294 & v4cb & v4cd & v5e & v406 & v4ce & v29d & v29f & v4cf & v30f & v4d0;
wire rnx2x69 = rnx2x68 || v4d1;
wire onx2x69 = onx2x68 || ( rnx2x68 && v4d1);
wire v4d2 = v38e == Advice_5;
wire v4d3 = Advice_2 == Advice_17;
wire v4d4 = v403 & v4d2 & v294 & v299 & v2d6 & v29f & v405 & v2f1 & v1e3 & v29d & v2e4 & v4d3;
wire rnx2x70 = rnx2x69 || v4d4;
wire onx2x70 = onx2x69 || ( rnx2x69 && v4d4);
wire v4d5 = v465 == Advice_5;
wire v4d6 = v4d5 & v403 & v299 & v2d6 & v406 & v294 & v1ef & v29d & v29f & v30f;
wire rnx2x71 = rnx2x70 || v4d6;
wire onx2x71 = onx2x70 || ( rnx2x70 && v4d6);
wire v4d7 = v4c0 == Advice_5;
wire v4d8 = v3a1 == Advice_21;
wire v4d9 = v3a1 == Advice_9;
wire v4da = Advice_9 == Advice_1;
wire [2:0] v4db = { Advice_21 , vd8 };
wire v4dc = v4db == Advice_14;
wire v4dd = v4ce & v4d7 & v294 & v2d6 & v299 & v4d8 & v29d & v4b6 & vd4 & v4d9 & v29f & v4da & v4b7 & v4dc;
wire rnx2x72 = rnx2x71 || v4dd;
wire onx2x72 = onx2x71 || ( rnx2x71 && v4dd);
wire v4de = v2ce & v245 & v248 & v2cf & v253 & v256 & v259 & v25c & v2da & v264 & v267 & v26a & v26d & v270 & v273 & v276 & v401 & v27e & v402 & v283 & v286 & v289;
wire [31:0] v4df = v4bd + v313;
wire [15:0] v4e0 = v4df[15:0];
wire [31:0] v4e1 = { 16'b0000000000000000, v4e0 };
wire v4e2 = v4e1 == Advice_5;
wire v4e3 = v4de & v2d6 & v4d8 & v4d9 & v4b6 & v4e2 & v294 & v299 & v17 & v29d & v29f & v4da & v4b7 & v4dc;
wire rnx2x73 = rnx2x72 || v4e3;
wire onx2x73 = onx2x72 || ( rnx2x72 && v4e3);
wire [31:0] v4e4 = v430 + v40f;
wire [31:0] v4e5 = v4e4 + v128;
wire v4e6 = v4e5 == Advice_5;
wire v4e7 = v40c == Advice_16;
wire v4e8 = v327 == Advice_3;
wire v4e9 = v40c == Advice_32;
wire v4ea = v294 & v299 & v297 & v2db & v4e6 & v4e7 & v201 & v4e8 & v4e9 & v29d & v29f & v4cf & v30f & v4d0;
wire rnx2x74 = rnx2x73 || v4ea;
wire onx2x74 = onx2x73 || ( rnx2x73 && v4ea);
wire v4eb = v35d == Advice_5;
wire v4ec = v2ec == Advice_2;
wire v4ed = v2b3 & v4eb & v294 & v299 & v4ec & v2ed & vef & v29d & v2b5 & v29f & v2e4 & v408;
wire rnx2x75 = rnx2x74 || v4ed;
wire onx2x75 = onx2x74 || ( rnx2x74 && v4ed);
wire v4ee = v352 == Advice_5;
wire v4ef = v2e9 & v299 & v2b5 & v4ec & v2ed & v4ee & v294 & v29f & vf8 & v29d & v2e4 & v408;
wire rnx2x76 = rnx2x75 || v4ef;
wire onx2x76 = onx2x75 || ( rnx2x75 && v4ef);
wire v4f0 = v44c == Advice_32;
wire [31:0] v4f1 = v431 + v30c;
wire v4f2 = v4f1 == Advice_5;
wire v4f3 = v44c == Advice_16;
wire v4f4 = v299 & v294 & v2b5 & v29d & v4f0 & v4f2 & v4f3 & v2f5 & ve9 & v29f & v4cf & v4d0;
wire rnx2x77 = rnx2x76 || v4f4;
wire onx2x77 = onx2x76 || ( rnx2x76 && v4f4);
wire v4f5 = v2a5 & v245 & v248 & v2a9 & v253 & v256 & v259 & v25c & v2da & v264 & v267 & v26a & v26d & v270 & v273 & v276 & v2b1 & v27e & v2b2 & v283 & v286 & v289;
wire [31:0] v4f6 = v350 + v378;
wire [31:0] v4f7 = v4f6 + v313;
wire v4f8 = v4f7 == Advice_5;
wire v4f9 = v37e == Advice_23;
wire v4fa = v4f5 & v4f8 & v294 & v405 & v2b5 & v4f9 & v299 & v2f1 & v29f & v1a4 & v29d & v2e4 & v3d5 & v408;
wire rnx2x78 = rnx2x77 || v4fa;
wire onx2x78 = onx2x77 || ( rnx2x77 && v4fa);
wire v4fb = v432 == Advice_5;
wire v4fc = v4fb & v2b5 & v4cb & v2f5 & v4cd & v294 & v18d & v299 & v29d & v29f & v4cf & v4d0;
wire rnx2x79 = rnx2x78 || v4fc;
wire onx2x79 = onx2x78 || ( rnx2x78 && v4fc);
wire v4fd = v387 == Advice_5;
wire v4fe = v4fd & v294 & v299 & v4f5 & v2b5 & v29d & v405 & v2f1 & vec & v29f & v2e4 & v408;
wire rnx2x80 = rnx2x79 || v4fe;
wire onx2x80 = onx2x79 || ( rnx2x79 && v4fe);
wire [31:0] v4ff = v3df + v28f;
wire v500 = v4ff == Advice_5;
wire v501 = v2a5 & v245 & v248 & v2a9 & v253 & v256 & v259 & v25c & v261 & v264 & v267 & v26a & v26d & v270 & v273 & v276 & v2b1 & v27e & v2b2 & v283 & v286 & v289;
wire v502 = v2e2 == Advice_2;
wire v503 = Advice_2 == Advice_24;
wire v504 = v294 & v500 & v299 & v501 & v502 & v4e8 & v2e3 & v2b5 & ve4 & v29d & v29f & v2e4 & v407 & v503;
wire rnx2x81 = rnx2x80 || v504;
wire onx2x81 = onx2x80 || ( rnx2x80 && v504);
wire v505 = v2a5 & v245 & v248 & v2a9 & v253 & v256 & v259 & v25c & v31f & v264 & v267 & v26a & v26d & v270 & v273 & v276 & v2b1 & v27e & v2b2 & v283 & v286 & v289;
wire v506 = v39f == Advice_5;
wire [2:0] v507 = { Advice_9 , vd8 };
wire v508 = v507 == Advice_18;
wire v509 = v294 & v4d8 & v299 & v4d9 & v4b6 & v505 & v506 & v2b5 & v14b & v29d & v29f & v508 & v4b7 & v4dc;
wire rnx2x82 = rnx2x81 || v509;
wire onx2x82 = onx2x81 || ( rnx2x81 && v509);
wire [31:0] v50a = v4a2 + v323;
wire v50b = v50a == Advice_5;
wire v50c = Advice_2 == Advice_31;
wire v50d = v505 & v299 & v294 & v502 & v29f & v4e8 & v50b & v2e3 & v2b5 & v13d & v29d & v2e4 & v407 & v50c;
wire rnx2x83 = rnx2x82 || v50d;
wire onx2x83 = onx2x82 || ( rnx2x82 && v50d);
wire v50e = v3ed == Advice_5;
wire v50f = Advice_9 == Advice_26;
wire [1:0] v510 = { Advice_21 , v11 };
wire v511 = v510 == Advice_25;
wire v512 = v294 & v299 & v2b5 & v4d8 & v50e & v4d9 & vf5 & v29d & v2f5 & v29f & v50f & v511;
wire rnx2x84 = rnx2x83 || v512;
wire onx2x84 = onx2x83 || ( rnx2x83 && v512);
wire [63:0] v513 = 64'b1111111111111111111111111111111100000000000000000000000000000000;
wire v514 = v23c > v513;
wire v515 = v514 == Out_register_CF;
wire v516 = v514 == Out_register_OF;
wire v517 = v2a5 & v245 & v248 & v2a9 & v253 & v256 & v259 & v25c & v2e8 & v264 & v267 & v26a & v26d & v270 & v273 & v276 & v515 & v27e & v516 & v283 & v286 & v289;
wire v518 = v517 & v2ea & v294 & v299 & v2ed & vcd & v29d & v29f & v2e4;
wire rnx2x85 = rnx2x84 || v518;
wire onx2x85 = onx2x84 || ( rnx2x84 && v518);
wire v519 = v2a5 & v245 & v248 & v2a9 & v253 & v256 & v259 & v25c & v2f4 & v264 & v267 & v26a & v26d & v270 & v273 & v276 & v515 & v27e & v516 & v283 & v286 & v289;
wire v51a = v294 & v29f & v299 & vc6 & v2ea & v2f1 & v519 & v29d & v2e4;
wire rnx2x86 = rnx2x85 || v51a;
wire onx2x86 = onx2x85 || ( rnx2x85 && v51a);
wire v51b = v2d4 & v4ec & v2ed & v4eb & v294 & v51 & v29d & v299 & v2d6 & v29f & v2e4 & v408;
wire rnx2x87 = rnx2x86 || v51b;
wire onx2x87 = onx2x86 || ( rnx2x86 && v51b);
wire v51c = v2ce & v245 & v248 & v2cf & v253 & v256 & v259 & v25c & v2f4 & v264 & v267 & v26a & v26d & v270 & v273 & v276 & v2d2 & v27e & v2d3 & v283 & v286 & v289;
wire [31:0] v51d = v4f6 + v128;
wire v51e = v51d == Advice_5;
wire v51f = v294 & v51c & v299 & v2d6 & v405 & v2f1 & v51e & v4f9 & v2d & v29d & v29f & v2e4 & v3d5 & v408;
wire rnx2x88 = rnx2x87 || v51f;
wire onx2x88 = onx2x87 || ( rnx2x87 && v51f);
wire v520 = v2ce & v245 & v248 & v2cf & v253 & v256 & v259 & v25c & v2b9 & v264 & v267 & v26a & v26d & v270 & v273 & v276 & v2d2 & v27e & v2d3 & v283 & v286 & v289;
wire [31:0] v521 = v4f6 + v2bb;
wire v522 = v521 == Advice_5;
wire v523 = v520 & v522 & v405 & v4f9 & v294 & v2d6 & v2f1 & v39 & v299 & v29d & v29f & v2e4 & v3d5 & v408;
wire rnx2x89 = rnx2x88 || v523;
wire onx2x89 = onx2x88 || ( rnx2x88 && v523);
wire v524 = v383 == Advice_5;
wire v525 = v520 & v524 & v299 & v2d6 & v405 & v2f1 & v294 & v29f & v9b & v29d & v2e4 & v408;
wire rnx2x90 = rnx2x89 || v525;
wire onx2x90 = onx2x89 || ( rnx2x89 && v525);
wire v526 = v520 & v4d5 & v2d6 & v1e9 & v299 & v406 & v29d & v294 & v29f & v30f;
wire rnx2x91 = rnx2x90 || v526;
wire onx2x91 = onx2x90 || ( rnx2x90 && v526);
wire v527 = v2ce & v245 & v248 & v2cf & v253 & v256 & v259 & v25c & v2da & v264 & v267 & v26a & v26d & v270 & v273 & v276 & v2d2 & v27e & v2d3 & v283 & v286 & v289;
wire v528 = v294 & v4e7 & v4e6 & v4e9 & v2d6 & v4e8 & v527 & v299 & v1d6 & v29d & v29f & v4cf & v30f & v4d0;
wire rnx2x92 = rnx2x91 || v528;
wire onx2x92 = onx2x91 || ( rnx2x91 && v528);
wire v529 = v519 & v4f2 & v299 & v4f3 & v4f0 & v1cf & v2b5 & v29d & v294 & v29f & v4cf & v4d0;
wire rnx2x93 = rnx2x92 || v529;
wire onx2x93 = onx2x92 || ( rnx2x92 && v529);
wire v52a = v517 & v4ee & v2b5 & v4ec & v299 & v29d & v2ed & v294 & v1cc & v29f & v2e4 & v408;
wire rnx2x94 = rnx2x93 || v52a;
wire onx2x94 = onx2x93 || ( rnx2x93 && v52a);
wire v52b = v373 == Advice_5;
wire v52c = v2a5 & v245 & v248 & v2a9 & v253 & v256 & v259 & v25c & v2da & v264 & v267 & v26a & v26d & v270 & v273 & v276 & v515 & v27e & v516 & v283 & v286 & v289;
wire v52d = v52b & v299 & v294 & v405 & v2b5 & v2f1 & v52c & v1bb & v406 & v29d & v29f & v2e4 & v407 & v408;
wire rnx2x95 = rnx2x94 || v52d;
wire onx2x95 = onx2x94 || ( rnx2x94 && v52d);
wire v52e = v519 & v294 & v2b5 & v405 & v4ee & v2f1 & v29f & v1c9 & v299 & v29d & v2e4 & v408;
wire rnx2x96 = rnx2x95 || v52e;
wire onx2x96 = onx2x95 || ( rnx2x95 && v52e);
wire v52f = v52c & v294 & v299 & v405 & v4fd & v2b5 & v1bc & v2f1 & v29d & v29f & v2e4 & v408;
wire rnx2x97 = rnx2x96 || v52f;
wire onx2x97 = onx2x96 || ( rnx2x96 && v52f);
wire v530 = v2a5 & v245 & v248 & v2a9 & v253 & v256 & v259 & v25c & v261 & v264 & v267 & v26a & v26d & v270 & v273 & v276 & v515 & v27e & v516 & v283 & v286 & v289;
wire v531 = v3bb == Advice_5;
wire v532 = v530 & v531 & v502 & v299 & v2e3 & v29f & v4e8 & v1bf & v294 & v2b5 & v29d & v2e4 & v407 & v4d3;
wire rnx2x98 = rnx2x97 || v532;
wire onx2x98 = onx2x97 || ( rnx2x97 && v532);
wire [31:0] v533 = v4c4 + v323;
wire v534 = v533 == Advice_5;
wire v535 = v2a5 & v245 & v248 & v2a9 & v253 & v256 & v259 & v25c & v31f & v264 & v267 & v26a & v26d & v270 & v273 & v276 & v515 & v27e & v516 & v283 & v286 & v289;
wire v536 = Advice_2 == Advice_30;
wire v537 = v534 & v299 & v535 & v502 & v294 & v2e3 & v29f & v1c2 & v4e8 & v2b5 & v29d & v2e4 & v407 & v536;
wire rnx2x99 = rnx2x98 || v537;
wire onx2x99 = onx2x98 || ( rnx2x98 && v537);
wire v2 = (!onx2x99) && rnx2x99;
assign result = v2;
assign dummy = 1'b0;
endmodule
